`timescale 1ns / 1ps
// A crude SRAM for testing with an initial state

module SRAM #(parameter ADR = 10, parameter DAT = 32, parameter DPTH = 1024)(
    output logic [DAT-1:0] DOUT,
    input logic [DAT-1:0] DIN,
    input logic [ADR-1:0] ADDR,
    input logic WE, RD, clk, rst_n
);
  
  //internal variables
  logic [DAT-1:0] SRAMs [DPTH-1:0];
  
  initial 
  begin
      //pre-load the image into SRAM
      $readmemh("image.txt", SRAMs);
  end

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      SRAMs[0]   <= 32'h21111111;
      SRAMs[1]   <= 32'h33322222;
      SRAMs[2]   <= 32'h44444333;
      SRAMs[3]   <= 32'h55555554;
      SRAMs[4]   <= 32'h77666666;
      SRAMs[5]   <= 32'h88887777;
      SRAMs[6]   <= 32'h99999988;
      SRAMs[7]   <= 32'hBAAAAAAA;
      SRAMs[8]   <= 32'h44141411;
      SRAMs[9]   <= 32'h44344424;
      SRAMs[10]  <= 32'h44444434;
      SRAMs[11]  <= 32'h44544454;
      SRAMs[12]  <= 32'h44744464;
      SRAMs[13]  <= 32'h88888774;
      SRAMs[14]  <= 32'h99999988;
      SRAMs[15]  <= 32'hBBAAAAAA;
      SRAMs[16]  <= 32'h00404041;
      SRAMs[17]  <= 32'h00400040;
      SRAMs[18]  <= 32'h00404040;
      SRAMs[19]  <= 32'h00400040;
      SRAMs[20]  <= 32'h00400040;
      SRAMs[21]  <= 32'h88888740;
      SRAMs[22]  <= 32'hA9999998;
      SRAMs[23]  <= 32'hBBAAAAAA;
      SRAMs[24]  <= 32'h40404041;
      SRAMs[25]  <= 32'h40440424;
      SRAMs[26]  <= 32'h04404044;
      SRAMs[27]  <= 32'h40404044;
      SRAMs[28]  <= 32'h40404464;
      SRAMs[29]  <= 32'h88888874;
      SRAMs[30]  <= 32'hA9999998;
      SRAMs[31]  <= 32'hBBBAAAAA;
      SRAMs[32]  <= 32'h00400041;
      SRAMs[33]  <= 32'h40440424;
      SRAMs[34]  <= 32'h04400043;
      SRAMs[35]  <= 32'h00400044;
      SRAMs[36]  <= 32'h00400040;
      SRAMs[37]  <= 32'h88888840;
      SRAMs[38]  <= 32'hAA999999;
      SRAMs[39]  <= 32'hBBBAAAAA;
      SRAMs[40]  <= 32'h40404041;
      SRAMs[41]  <= 32'h40440424;
      SRAMs[42]  <= 32'h04404044;
      SRAMs[43]  <= 32'h44644044;
      SRAMs[44]  <= 32'h44744040;
      SRAMs[45]  <= 32'h88888840;
      SRAMs[46]  <= 32'hAA999999;
      SRAMs[47]  <= 32'hBBBBAAAA;
      SRAMs[48]  <= 32'h00404041;
      SRAMs[49]  <= 32'h00400040;
      SRAMs[50]  <= 32'h00404040;
      SRAMs[51]  <= 32'h00454040;
      SRAMs[52]  <= 32'h00400040;
      SRAMs[53]  <= 32'h98888840;
      SRAMs[54]  <= 32'hAAA99999;
      SRAMs[55]  <= 32'hBBBBAAAA;
      SRAMs[56]  <= 32'h44242411;
      SRAMs[57]  <= 32'h44344434;
      SRAMs[58]  <= 32'h44444444;
      SRAMs[59]  <= 32'h44665454;
      SRAMs[60]  <= 32'h44744464;
      SRAMs[61]  <= 32'h98888884;
      SRAMs[62]  <= 32'hAAA99999;
      SRAMs[63]  <= 32'hBBBBBAAA;
      SRAMs[64]  <= 32'h22222111;
      SRAMs[65]  <= 32'h43333332;
      SRAMs[66]  <= 32'h55544444;
      SRAMs[67]  <= 32'h66665555;
      SRAMs[68]  <= 32'h77777766;
      SRAMs[69]  <= 32'h99888888;
      SRAMs[70]  <= 32'hAAAA9999;
      SRAMs[71]  <= 32'hBBBBBAAA;
      SRAMs[72]  <= 32'h22222211;
      SRAMs[73]  <= 32'h43333333;
      SRAMs[74]  <= 32'h55544444;
      SRAMs[75]  <= 32'h66666555;
      SRAMs[76]  <= 32'h87777776;
      SRAMs[77]  <= 32'h99888888;
      SRAMs[78]  <= 32'hAAAA9999;
      SRAMs[79]  <= 32'hBBBBBBAA;
      SRAMs[80]  <= 32'h22222211;
      SRAMs[81]  <= 32'h44333333;
      SRAMs[82]  <= 32'h55554444;
      SRAMs[83]  <= 32'h66666555;
      SRAMs[84]  <= 32'h87777776;
      SRAMs[85]  <= 32'h99988888;
      SRAMs[86]  <= 32'hAAAAA999;
      SRAMs[87]  <= 32'hBBBBBBAA;
      SRAMs[88]  <= 32'h32222221;
      SRAMs[89]  <= 32'h44333333;
      SRAMs[90]  <= 32'h55554444;
      SRAMs[91]  <= 32'h66666655;
      SRAMs[92]  <= 32'h88777777;
      SRAMs[93]  <= 32'h99988888;
      SRAMs[94]  <= 32'hAAAAA999;
      SRAMs[95]  <= 32'hCBBBBBBA;
      SRAMs[96]  <= 32'h32222221;
      SRAMs[97]  <= 32'h44433333;
      SRAMs[98]  <= 32'h55555444;
      SRAMs[99]  <= 32'h66666655;
      SRAMs[100] <= 32'h88777777;
      SRAMs[101] <= 32'h99998888;
      SRAMs[102] <= 32'hAAAAAA99;
      SRAMs[103] <= 32'hCBBBBBBA;
      SRAMs[104] <= 32'h33222222;
      SRAMs[105] <= 32'h44433333;
      SRAMs[106] <= 32'h55555444;
      SRAMs[107] <= 32'h76666665;
      SRAMs[108] <= 32'h88877777;
      SRAMs[109] <= 32'h99998888;
      SRAMs[110] <= 32'hAAAAAA99;
      SRAMs[111] <= 32'hCCBBBBBB;
      SRAMs[112] <= 32'h33222222;
      SRAMs[113] <= 32'h44443333;
      SRAMs[114] <= 32'h55555544;
      SRAMs[115] <= 32'h76666665;
      SRAMs[116] <= 32'h88877777;
      SRAMs[117] <= 32'h99999888;
      SRAMs[118] <= 32'hAAAAAAA9;
      SRAMs[119] <= 32'hCCBBBBBB;
      SRAMs[120] <= 32'h33322222;
      SRAMs[121] <= 32'h44443333;
      SRAMs[122] <= 32'h55555544;
      SRAMs[123] <= 32'h77666666;
      SRAMs[124] <= 32'h88887777;
      SRAMs[125] <= 32'h99999888;
      SRAMs[126] <= 32'hBAAAAAA9;
      SRAMs[127] <= 32'hCCCBBBBB;
      SRAMs[128] <= 32'h33322222;
      SRAMs[129] <= 32'h44444333;
      SRAMs[130] <= 32'h55555554;
      SRAMs[131] <= 32'h77666666;
      SRAMs[132] <= 32'h88887777;
      SRAMs[133] <= 32'h99999988;
      SRAMs[134] <= 32'hBAAAAAAA;
      SRAMs[135] <= 32'hCCCBBBBB;
      SRAMs[136] <= 32'h33332222;
      SRAMs[137] <= 32'h44444333;
      SRAMs[138] <= 32'h65555554;
      SRAMs[139] <= 32'h77766666;
      SRAMs[140] <= 32'h88888777;
      SRAMs[141] <= 32'h99999988;
      SRAMs[142] <= 32'hBBAAAAAA;
      SRAMs[143] <= 32'hCCCCBBBB;
      SRAMs[144] <= 32'h33332222;
      SRAMs[145] <= 32'h44444433;
      SRAMs[146] <= 32'h65555555;
      SRAMs[147] <= 32'h77766666;
      SRAMs[148] <= 32'h88888777;
      SRAMs[149] <= 32'hA9999998;
      SRAMs[150] <= 32'hBBAAAAAA;
      SRAMs[151] <= 32'hCCCCBBBB;
      SRAMs[152] <= 32'h55353522;
      SRAMs[153] <= 32'h55455535;
      SRAMs[154] <= 32'h65555555;
      SRAMs[155] <= 32'h55775566;
      SRAMs[156] <= 32'h55855575;
      SRAMs[157] <= 32'hA9999995;
      SRAMs[158] <= 32'hBBBAAAAA;
      SRAMs[159] <= 32'hCCCCCBBB;
      SRAMs[160] <= 32'h00505052;
      SRAMs[161] <= 32'h00500050;
      SRAMs[162] <= 32'h50500055;
      SRAMs[163] <= 32'h00550056;
      SRAMs[164] <= 32'h00500050;
      SRAMs[165] <= 32'hAA999950;
      SRAMs[166] <= 32'hBBBAAAAA;
      SRAMs[167] <= 32'hCCCCCBBB;
      SRAMs[168] <= 32'h50505052;
      SRAMs[169] <= 32'h50550545;
      SRAMs[170] <= 32'h50555050;
      SRAMs[171] <= 32'h50505056;
      SRAMs[172] <= 32'h50505055;
      SRAMs[173] <= 32'hAA999995;
      SRAMs[174] <= 32'hBBBBAAAA;
      SRAMs[175] <= 32'hCCCCCCBB;
      SRAMs[176] <= 32'h00500052;
      SRAMs[177] <= 32'h50550545;
      SRAMs[178] <= 32'h50550050;
      SRAMs[179] <= 32'h00550056;
      SRAMs[180] <= 32'h50500055;
      SRAMs[181] <= 32'hAAA99950;
      SRAMs[182] <= 32'hBBBBAAAA;
      SRAMs[183] <= 32'hCCCCCCBB;
      SRAMs[184] <= 32'h50505052;
      SRAMs[185] <= 32'h50550545;
      SRAMs[186] <= 32'h50555050;
      SRAMs[187] <= 32'h50505055;
      SRAMs[188] <= 32'h50550055;
      SRAMs[189] <= 32'hAAA99950;
      SRAMs[190] <= 32'hBBBBBAAA;
      SRAMs[191] <= 32'hCCCCCCCB;
      SRAMs[192] <= 32'h00505052;
      SRAMs[193] <= 32'h00500050;
      SRAMs[194] <= 32'h00500055;
      SRAMs[195] <= 32'h00550050;
      SRAMs[196] <= 32'h00505050;
      SRAMs[197] <= 32'hAAAA9950;
      SRAMs[198] <= 32'hBBBBBAAA;
      SRAMs[199] <= 32'hDCCCCCCB;
      SRAMs[200] <= 32'h55353533;
      SRAMs[201] <= 32'h55555545;
      SRAMs[202] <= 32'h55655555;
      SRAMs[203] <= 32'h55775575;
      SRAMs[204] <= 32'h55858585;
      SRAMs[205] <= 32'hAAAA9995;
      SRAMs[206] <= 32'hBBBBBBAA;
      SRAMs[207] <= 32'hDCCCCCCC;
      SRAMs[208] <= 32'h44333333;
      SRAMs[209] <= 32'h55554444;
      SRAMs[210] <= 32'h66666555;
      SRAMs[211] <= 32'h87777776;
      SRAMs[212] <= 32'h99988888;
      SRAMs[213] <= 32'hAAAAA999;
      SRAMs[214] <= 32'hBBBBBBAA;
      SRAMs[215] <= 32'hDDCCCCCC;
      SRAMs[216] <= 32'h44333333;
      SRAMs[217] <= 32'h55554444;
      SRAMs[218] <= 32'h66666655;
      SRAMs[219] <= 32'h88777777;
      SRAMs[220] <= 32'h99988888;
      SRAMs[221] <= 32'hAAAAA999;
      SRAMs[222] <= 32'hCBBBBBBA;
      SRAMs[223] <= 32'hDDCCCCCC;
      SRAMs[224] <= 32'h44433333;
      SRAMs[225] <= 32'h55555444;
      SRAMs[226] <= 32'h66666655;
      SRAMs[227] <= 32'h88777777;
      SRAMs[228] <= 32'h99998888;
      SRAMs[229] <= 32'hAAAAAA99;
      SRAMs[230] <= 32'hCBBBBBBA;
      SRAMs[231] <= 32'hDDDCCCCC;
      SRAMs[232] <= 32'h44433333;
      SRAMs[233] <= 32'h55555444;
      SRAMs[234] <= 32'h76666665;
      SRAMs[235] <= 32'h88877777;
      SRAMs[236] <= 32'h99998888;
      SRAMs[237] <= 32'hAAAAAA99;
      SRAMs[238] <= 32'hCCBBBBBB;
      SRAMs[239] <= 32'hDDDCCCCC;
      SRAMs[240] <= 32'h44443333;
      SRAMs[241] <= 32'h55555544;
      SRAMs[242] <= 32'h76666665;
      SRAMs[243] <= 32'h88877777;
      SRAMs[244] <= 32'h99999888;
      SRAMs[245] <= 32'hAAAAAAA9;
      SRAMs[246] <= 32'hCCBBBBBB;
      SRAMs[247] <= 32'hDDDDCCCC;
      SRAMs[248] <= 32'h44443333;
      SRAMs[249] <= 32'h55555544;
      SRAMs[250] <= 32'h77666666;
      SRAMs[251] <= 32'h88887777;
      SRAMs[252] <= 32'h99999888;
      SRAMs[253] <= 32'hBAAAAAA9;
      SRAMs[254] <= 32'hCCCBBBBB;
      SRAMs[255] <= 32'hDDDDCCCC;
      SRAMs[256] <= 32'h44444333;
      SRAMs[257] <= 32'h55555554;
      SRAMs[258] <= 32'h77666666;
      SRAMs[259] <= 32'h88887777;
      SRAMs[260] <= 32'h99999988;
      SRAMs[261] <= 32'hBAAAAAAA;
      SRAMs[262] <= 32'hCCCBBBBB;
      SRAMs[263] <= 32'hDDDDDCCC;
      SRAMs[264] <= 32'h44422233;
      SRAMs[265] <= 32'h65522254;
      SRAMs[266] <= 32'h72722266;
      SRAMs[267] <= 32'h88822272;
      SRAMs[268] <= 32'h22922288;
      SRAMs[269] <= 32'hBBAAAAA2;
      SRAMs[270] <= 32'hCCCCBBBB;
      SRAMs[271] <= 32'hDDDDDCCC;
      SRAMs[272] <= 32'h44200023;
      SRAMs[273] <= 32'h65200025;
      SRAMs[274] <= 32'h20200026;
      SRAMs[275] <= 32'h88200020;
      SRAMs[276] <= 32'h00200028;
      SRAMs[277] <= 32'hBBAAAA20;
      SRAMs[278] <= 32'hCCCCBBBB;
      SRAMs[279] <= 32'hDDDDDDCC;
      SRAMs[280] <= 32'h22202233;
      SRAMs[281] <= 32'h66202022;
      SRAMs[282] <= 32'h20202026;
      SRAMs[283] <= 32'h88822020;
      SRAMs[284] <= 32'h20202298;
      SRAMs[285] <= 32'hBBBAAAA2;
      SRAMs[286] <= 32'hCCCCCBBB;
      SRAMs[287] <= 32'hDDDDDDCC;
      SRAMs[288] <= 32'h00200023;
      SRAMs[289] <= 32'h66200020;
      SRAMs[290] <= 32'h20200026;
      SRAMs[291] <= 32'h88202020;
      SRAMs[292] <= 32'h00200029;
      SRAMs[293] <= 32'hBBBAAA20;
      SRAMs[294] <= 32'hCCCCCBBB;
      SRAMs[295] <= 32'hEDDDDDDC;
      SRAMs[296] <= 32'h22202243;
      SRAMs[297] <= 32'h66202022;
      SRAMs[298] <= 32'h20202026;
      SRAMs[299] <= 32'h88202020;
      SRAMs[300] <= 32'h22922029;
      SRAMs[301] <= 32'hBBBBAA20;
      SRAMs[302] <= 32'hCCCCCCBB;
      SRAMs[303] <= 32'hEDDDDDDC;
      SRAMs[304] <= 32'h55200024;
      SRAMs[305] <= 32'h66200025;
      SRAMs[306] <= 32'h00202026;
      SRAMs[307] <= 32'h98200020;
      SRAMs[308] <= 32'h00200029;
      SRAMs[309] <= 32'hBBBBAA20;
      SRAMs[310] <= 32'hCCCCCCBB;
      SRAMs[311] <= 32'hEEDDDDDD;
      SRAMs[312] <= 32'h55422244;
      SRAMs[313] <= 32'h66622255;
      SRAMs[314] <= 32'h22727266;
      SRAMs[315] <= 32'h98822282;
      SRAMs[316] <= 32'h22A22299;
      SRAMs[317] <= 32'hBBBBBAA2;
      SRAMs[318] <= 32'hCCCCCCCB;
      SRAMs[319] <= 32'hEEDDDDDD;
      SRAMs[320] <= 32'h55544444;
      SRAMs[321] <= 32'h66665555;
      SRAMs[322] <= 32'h77777766;
      SRAMs[323] <= 32'h99888888;
      SRAMs[324] <= 32'hAAAA9999;
      SRAMs[325] <= 32'hBBBBBAAA;
      SRAMs[326] <= 32'hDCCCCCCB;
      SRAMs[327] <= 32'hEEEDDDDD;
      SRAMs[328] <= 32'h55544444;
      SRAMs[329] <= 32'h66666555;
      SRAMs[330] <= 32'h87777776;
      SRAMs[331] <= 32'h99888888;
      SRAMs[332] <= 32'hAAAA9999;
      SRAMs[333] <= 32'hBBBBBBAA;
      SRAMs[334] <= 32'hDCCCCCCC;
      SRAMs[335] <= 32'hEEEDDDDD;
      SRAMs[336] <= 32'h55554444;
      SRAMs[337] <= 32'h66666555;
      SRAMs[338] <= 32'h87777776;
      SRAMs[339] <= 32'h99988888;
      SRAMs[340] <= 32'hAAAAA999;
      SRAMs[341] <= 32'hBBBBBBAA;
      SRAMs[342] <= 32'hDDCCCCCC;
      SRAMs[343] <= 32'hEEEEDDDD;
      SRAMs[344] <= 32'h55554444;
      SRAMs[345] <= 32'h66666655;
      SRAMs[346] <= 32'h88777777;
      SRAMs[347] <= 32'h99988888;
      SRAMs[348] <= 32'hAAAAA999;
      SRAMs[349] <= 32'hCBBBBBBA;
      SRAMs[350] <= 32'hDDCCCCCC;
      SRAMs[351] <= 32'hEEEEDDDD;
      SRAMs[352] <= 32'h55555444;
      SRAMs[353] <= 32'h66666655;
      SRAMs[354] <= 32'h88777777;
      SRAMs[355] <= 32'h99998888;
      SRAMs[356] <= 32'hAAAAAA99;
      SRAMs[357] <= 32'hCBBBBBBA;
      SRAMs[358] <= 32'hDDDCCCCC;
      SRAMs[359] <= 32'hEEEEEDDD;
      SRAMs[360] <= 32'h55555444;
      SRAMs[361] <= 32'h76666665;
      SRAMs[362] <= 32'h88877777;
      SRAMs[363] <= 32'h99998888;
      SRAMs[364] <= 32'hAAAAAA99;
      SRAMs[365] <= 32'hCCBBBBBB;
      SRAMs[366] <= 32'hDDDCCCCC;
      SRAMs[367] <= 32'hEEEEEDDD;
      SRAMs[368] <= 32'h55555544;
      SRAMs[369] <= 32'h76666665;
      SRAMs[370] <= 32'h88877777;
      SRAMs[371] <= 32'h99999888;
      SRAMs[372] <= 32'hAAAAAAA9;
      SRAMs[373] <= 32'hCCBBBBBB;
      SRAMs[374] <= 32'hDDDDCCCC;
      SRAMs[375] <= 32'hEEEEEEDD;
      SRAMs[376] <= 32'h55555544;
      SRAMs[377] <= 32'h77666666;
      SRAMs[378] <= 32'h88887777;
      SRAMs[379] <= 32'h99999888;
      SRAMs[380] <= 32'hBAAAAAA9;
      SRAMs[381] <= 32'hCCCBBBBB;
      SRAMs[382] <= 32'hDDDDCCCC;
      SRAMs[383] <= 32'hEEEEEEDD;
      
      //SRAMs[0:383] <= {32'h11111112, 32'h22222333, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'h11414144, 32'h42444344, 32'h43444444, 32'h45444544, 32'h46444777, 32'h77788888, 32'h88999999, 32'hAAAAAABB, 32'h14040400, 32'h04000400, 32'h04040400, 32'h04000400, 32'h04000477, 32'h77788888, 32'h8999999A, 32'hAAAAAABB, 32'h14040404, 32'h42404404, 32'h44040440, 32'h44040404, 32'h46440477, 32'h77888888, 32'h8999999A, 32'hAAAAABBB, 32'h14000400, 32'h42404404, 32'h34000440, 32'h44000400, 32'h04000477, 32'h77888888, 32'h999999AA, 32'hAAAAABBB, 32'h14040404, 32'h42404404, 32'h44040440, 32'h44044644, 32'h04044777, 32'h78888888, 32'h999999AA, 32'hAAAABBBB, 32'h14040400, 32'h04000400, 32'h04040400, 32'h04045400, 32'h04000477, 32'h78888889, 32'h99999AAA, 32'hAAAABBBB, 32'h11424244, 32'h43444344, 32'h44444444, 32'h45456644, 32'h46444777, 32'h88888889, 32'h99999AAA, 32'hAAABBBBB, 32'h11122222, 32'h23333334, 32'h44444555, 32'h55556666, 32'h66777777, 32'h88888899, 32'h9999AAAA, 32'hAAABBBBB, 32'h11222222, 32'h33333334, 32'h44444555, 32'h55566666, 32'h67777778, 32'h88888899, 32'h9999AAAA, 32'hAABBBBBB, 32'h11222222, 32'h33333344, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'h12222223, 32'h33333344, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'h12222223, 32'h33333444, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'h22222233, 32'h33333444, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'h22222233, 32'h33334444, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'h22222333, 32'h33334444, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'h22222333, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'hBBBBBCCC, 32'h22223333, 32'h33344444, 32'h45555556, 32'h66666777, 32'h77788888, 32'h88999999, 32'hAAAAAABB, 32'hBBBBCCCC, 32'h22223333, 32'h33444444, 32'h55555556, 32'h66666777, 32'h77788888, 32'h8999999A, 32'hAAAAAABB, 32'hBBBBCCCC, 32'h22535355, 32'h53555455, 32'h55555556, 32'h66557755, 32'h57555855, 32'h5999999A, 32'hAAAAABBB, 32'hBBBCCCCC, 32'h25050500, 32'h05000500, 32'h55000505, 32'h65005500, 32'h05000500, 32'h059999AA, 32'hAAAAABBB, 32'hBBBCCCCC, 32'h25050505, 32'h54505505, 32'h05055505, 32'h65050505, 32'h55050505, 32'h599999AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'h25000500, 32'h54505505, 32'h05005505, 32'h65005500, 32'h55000505, 32'h05999AAA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'h25050505, 32'h54505505, 32'h05055505, 32'h55050505, 32'h55005505, 32'h05999AAA, 32'hAAABBBBB, 32'hBCCCCCCC, 32'h25050500, 32'h05000500, 32'h55000500, 32'h05005500, 32'h05050500, 32'h0599AAAA, 32'hAAABBBBB, 32'hBCCCCCCD, 32'h33535355, 32'h54555555, 32'h55555655, 32'h57557755, 32'h58585855, 32'h5999AAAA, 32'hAABBBBBB, 32'hCCCCCCCD, 32'h33333344, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'hCCCCCCDD, 32'h33333344, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'hCCCCCCDD, 32'h33333444, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'hCCCCCDDD, 32'h33333444, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'hCCCCCDDD, 32'h33334444, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'hCCCCDDDD, 32'h33334444, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'hCCCCDDDD, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'hBBBBBCCC, 32'hCCCDDDDD, 32'h33222444, 32'h45222556, 32'h66222727, 32'h27222888, 32'h88222999, 32'hAAAAAABB, 32'hBBBBCCCC, 32'hCCCDDDDD, 32'h32000244, 32'h52000256, 32'h62000202, 32'h02000288, 32'h8200029A, 32'hAAAAAABB, 32'hBBBBCCCC, 32'hCCDDDDDD, 32'h33220222, 32'h22020266, 32'h62020202, 32'h02022888, 32'h8922029A, 32'hAAAAABBB, 32'hBBBCCCCC, 32'hCCDDDDDD, 32'h32000200, 32'h02000266, 32'h62000202, 32'h02020288, 32'h920002AA, 32'hAAAAABBB, 32'hBBBCCCCC, 32'hCDDDDDDE, 32'h34220222, 32'h22020266, 32'h62020202, 32'h02020288, 32'h920229AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'hCDDDDDDE, 32'h42000255, 32'h52000266, 32'h62020200, 32'h02000289, 32'h920002AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'hDDDDDDEE, 32'h44222455, 32'h55222666, 32'h66272722, 32'h28222889, 32'h99222AAA, 32'hAAABBBBB, 32'hBCCCCCCC, 32'hDDDDDDEE, 32'h44444555, 32'h55556666, 32'h66777777, 32'h88888899, 32'h9999AAAA, 32'hAAABBBBB, 32'hBCCCCCCD, 32'hDDDDDEEE, 32'h44444555, 32'h55566666, 32'h67777778, 32'h88888899, 32'h9999AAAA, 32'hAABBBBBB, 32'hCCCCCCCD, 32'hDDDDDEEE, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'hCCCCCCDD, 32'hDDDDEEEE, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'hCCCCCCDD, 32'hDDDDEEEE, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'hCCCCCDDD, 32'hDDDEEEEE, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'hCCCCCDDD, 32'hDDDEEEEE, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'hCCCCDDDD, 32'hDDEEEEEE, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'hCCCCDDDD, 32'hDDEEEEEE};
    end
    else if (WE == 1'b1 && RD == 1'b0) SRAMs[ADDR] <= DIN;
    else;
  end

  assign DOUT = SRAMs[ADDR];

endmodule
