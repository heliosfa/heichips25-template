module heichips25_bagel (clk,
    ena,
    rst_n,
    tmds_b,
    tmds_clk,
    tmds_g,
    tmds_r,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 output tmds_b;
 output tmds_clk;
 output tmds_g;
 output tmds_r;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire clk_regs;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire \blue_tmds_par[0] ;
 wire \blue_tmds_par[1] ;
 wire \blue_tmds_par[2] ;
 wire \blue_tmds_par[3] ;
 wire \blue_tmds_par[5] ;
 wire \blue_tmds_par[6] ;
 wire \blue_tmds_par[7] ;
 wire \blue_tmds_par[8] ;
 wire \blue_tmds_par[9] ;
 wire clk_video;
 wire \clockdiv.q0 ;
 wire \clockdiv.q1 ;
 wire \clockdiv.q2 ;
 wire \clockdiv.q2temp ;
 wire display_enable;
 wire \green_tmds_par[0] ;
 wire \green_tmds_par[1] ;
 wire \green_tmds_par[2] ;
 wire \green_tmds_par[6] ;
 wire \green_tmds_par[7] ;
 wire \green_tmds_par[8] ;
 wire \green_tmds_par[9] ;
 wire hsync;
 wire \red_tmds_par[0] ;
 wire \red_tmds_par[1] ;
 wire \red_tmds_par[2] ;
 wire \red_tmds_par[3] ;
 wire \red_tmds_par[4] ;
 wire \red_tmds_par[5] ;
 wire \red_tmds_par[6] ;
 wire \red_tmds_par[7] ;
 wire \red_tmds_par[8] ;
 wire \red_tmds_par[9] ;
 wire \serialize.bit_cnt[0] ;
 wire \serialize.bit_cnt[1] ;
 wire \serialize.n410 ;
 wire \serialize.n411[0] ;
 wire \serialize.n411[1] ;
 wire \serialize.n411[2] ;
 wire \serialize.n411[3] ;
 wire \serialize.n411[4] ;
 wire \serialize.n411[5] ;
 wire \serialize.n411[6] ;
 wire \serialize.n411[7] ;
 wire \serialize.n414[0] ;
 wire \serialize.n414[1] ;
 wire \serialize.n414[2] ;
 wire \serialize.n414[3] ;
 wire \serialize.n414[4] ;
 wire \serialize.n414[5] ;
 wire \serialize.n414[6] ;
 wire \serialize.n414[7] ;
 wire \serialize.n417[0] ;
 wire \serialize.n417[1] ;
 wire \serialize.n417[2] ;
 wire \serialize.n417[3] ;
 wire \serialize.n417[4] ;
 wire \serialize.n417[5] ;
 wire \serialize.n417[6] ;
 wire \serialize.n417[7] ;
 wire \serialize.n420[0] ;
 wire \serialize.n420[1] ;
 wire \serialize.n420[2] ;
 wire \serialize.n420[3] ;
 wire \serialize.n420[4] ;
 wire \serialize.n420[6] ;
 wire \serialize.n427[0] ;
 wire \serialize.n427[1] ;
 wire \serialize.n427[2] ;
 wire \serialize.n427[3] ;
 wire \serialize.n427[4] ;
 wire \serialize.n427[5] ;
 wire \serialize.n427[6] ;
 wire \serialize.n427[7] ;
 wire \serialize.n427[8] ;
 wire \serialize.n427[9] ;
 wire \serialize.n428[0] ;
 wire \serialize.n428[1] ;
 wire \serialize.n428[2] ;
 wire \serialize.n428[3] ;
 wire \serialize.n428[4] ;
 wire \serialize.n428[5] ;
 wire \serialize.n428[6] ;
 wire \serialize.n428[7] ;
 wire \serialize.n428[8] ;
 wire \serialize.n428[9] ;
 wire \serialize.n429[0] ;
 wire \serialize.n429[1] ;
 wire \serialize.n429[2] ;
 wire \serialize.n429[3] ;
 wire \serialize.n429[4] ;
 wire \serialize.n429[5] ;
 wire \serialize.n429[6] ;
 wire \serialize.n429[7] ;
 wire \serialize.n429[8] ;
 wire \serialize.n429[9] ;
 wire \serialize.n431[0] ;
 wire \serialize.n431[1] ;
 wire \serialize.n431[2] ;
 wire \serialize.n431[3] ;
 wire \serialize.n431[4] ;
 wire \serialize.n431[5] ;
 wire \serialize.n431[6] ;
 wire \serialize.n433[0] ;
 wire \serialize.n433[1] ;
 wire \serialize.n450 ;
 wire \serialize.n452 ;
 wire \serialize.n453 ;
 wire \serialize.n455 ;
 wire \serialize.n456 ;
 wire \serialize.n458 ;
 wire \serialize.n459 ;
 wire \serialize.n461 ;
 wire net3;
 wire \tmds_blue.dc_balancing_reg[0] ;
 wire \tmds_blue.dc_balancing_reg[1] ;
 wire \tmds_blue.dc_balancing_reg[2] ;
 wire \tmds_blue.dc_balancing_reg[3] ;
 wire \tmds_blue.dc_balancing_reg[4] ;
 wire \tmds_blue.n100 ;
 wire \tmds_blue.n126 ;
 wire \tmds_blue.n132 ;
 wire \tmds_blue.n193 ;
 wire \tmds_blue.vsync ;
 wire net4;
 wire net5;
 wire \tmds_green.dc_balancing_reg[0] ;
 wire \tmds_green.dc_balancing_reg[1] ;
 wire \tmds_green.dc_balancing_reg[2] ;
 wire \tmds_green.dc_balancing_reg[3] ;
 wire \tmds_green.dc_balancing_reg[4] ;
 wire \tmds_green.n100 ;
 wire \tmds_green.n126 ;
 wire \tmds_green.n132 ;
 wire net6;
 wire \tmds_red.dc_balancing_reg[0] ;
 wire \tmds_red.dc_balancing_reg[1] ;
 wire \tmds_red.dc_balancing_reg[2] ;
 wire \tmds_red.dc_balancing_reg[3] ;
 wire \tmds_red.dc_balancing_reg[4] ;
 wire \tmds_red.n100 ;
 wire \tmds_red.n102 ;
 wire \tmds_red.n114 ;
 wire \tmds_red.n126 ;
 wire \tmds_red.n132 ;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net7;
 wire net30;
 wire net8;
 wire net9;
 wire net10;
 wire net31;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire \videogen.fancy_shader.n646[0] ;
 wire \videogen.fancy_shader.n646[1] ;
 wire \videogen.fancy_shader.n646[2] ;
 wire \videogen.fancy_shader.n646[3] ;
 wire \videogen.fancy_shader.n646[4] ;
 wire \videogen.fancy_shader.n646[5] ;
 wire \videogen.fancy_shader.n646[6] ;
 wire \videogen.fancy_shader.n646[7] ;
 wire \videogen.fancy_shader.n646[8] ;
 wire \videogen.fancy_shader.n646[9] ;
 wire \videogen.fancy_shader.video_x[0] ;
 wire \videogen.fancy_shader.video_x[1] ;
 wire \videogen.fancy_shader.video_x[2] ;
 wire \videogen.fancy_shader.video_x[3] ;
 wire \videogen.fancy_shader.video_x[4] ;
 wire \videogen.fancy_shader.video_x[5] ;
 wire \videogen.fancy_shader.video_x[6] ;
 wire \videogen.fancy_shader.video_x[7] ;
 wire \videogen.fancy_shader.video_x[8] ;
 wire \videogen.fancy_shader.video_x[9] ;
 wire \videogen.fancy_shader.video_y[0] ;
 wire \videogen.fancy_shader.video_y[1] ;
 wire \videogen.fancy_shader.video_y[2] ;
 wire \videogen.fancy_shader.video_y[3] ;
 wire \videogen.fancy_shader.video_y[4] ;
 wire \videogen.fancy_shader.video_y[5] ;
 wire \videogen.fancy_shader.video_y[6] ;
 wire \videogen.fancy_shader.video_y[7] ;
 wire \videogen.fancy_shader.video_y[8] ;
 wire \videogen.fancy_shader.video_y[9] ;
 wire \videogen.mem_read ;
 wire \videogen.mem_row ;
 wire \videogen.test_lut_thingy.gol_counter_reg[0] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[1] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[2] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net1;
 wire net2;
 wire net21;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;

 sg13g2_inv_1 _2514_ (.Y(_0632_),
    .A(\videogen.fancy_shader.video_y[9] ));
 sg13g2_inv_1 _2515_ (.Y(_0633_),
    .A(\videogen.fancy_shader.video_y[5] ));
 sg13g2_inv_1 _2516_ (.Y(_0634_),
    .A(\videogen.fancy_shader.n646[5] ));
 sg13g2_inv_1 _2517_ (.Y(_0635_),
    .A(\videogen.fancy_shader.n646[0] ));
 sg13g2_inv_4 _2518_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .Y(_0636_));
 sg13g2_inv_2 _2519_ (.Y(_0637_),
    .A(net612));
 sg13g2_inv_1 _2520_ (.Y(_0638_),
    .A(net614));
 sg13g2_inv_1 _2521_ (.Y(_0639_),
    .A(net619));
 sg13g2_inv_1 _2522_ (.Y(_0640_),
    .A(\videogen.fancy_shader.video_x[5] ));
 sg13g2_inv_1 _2523_ (.Y(_0641_),
    .A(\tmds_green.dc_balancing_reg[3] ));
 sg13g2_inv_2 _2524_ (.Y(_0642_),
    .A(\tmds_green.dc_balancing_reg[4] ));
 sg13g2_inv_2 _2525_ (.Y(_0643_),
    .A(net604));
 sg13g2_inv_1 _2526_ (.Y(_0644_),
    .A(\tmds_blue.dc_balancing_reg[4] ));
 sg13g2_inv_1 _2527_ (.Y(_0645_),
    .A(\tmds_blue.dc_balancing_reg[1] ));
 sg13g2_inv_1 _2528_ (.Y(_0646_),
    .A(\tmds_blue.dc_balancing_reg[3] ));
 sg13g2_inv_4 _2529_ (.A(net606),
    .Y(_0647_));
 sg13g2_inv_2 _2530_ (.Y(_0648_),
    .A(net793));
 sg13g2_inv_8 _2531_ (.Y(_0649_),
    .A(net600));
 sg13g2_inv_1 _2532_ (.Y(_0650_),
    .A(net2));
 sg13g2_inv_1 _2533_ (.Y(_0651_),
    .A(\videogen.test_lut_thingy.gol_counter_reg[2] ));
 sg13g2_inv_1 _2534_ (.Y(_0652_),
    .A(\tmds_red.dc_balancing_reg[4] ));
 sg13g2_inv_1 _2535_ (.Y(_0653_),
    .A(\tmds_red.dc_balancing_reg[3] ));
 sg13g2_inv_1 _2536_ (.Y(_0654_),
    .A(\tmds_red.dc_balancing_reg[2] ));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_inv_1 _2538_ (.Y(_0655_),
    .A(net417));
 sg13g2_inv_1 _2539_ (.Y(_0656_),
    .A(net414));
 sg13g2_inv_1 _2540_ (.Y(_0657_),
    .A(net421));
 sg13g2_nand2_1 _2541_ (.Y(_0658_),
    .A(net429),
    .B(net413));
 sg13g2_xor2_1 _2542_ (.B(net413),
    .A(net429),
    .X(\serialize.n433[1] ));
 sg13g2_nand2_1 _2543_ (.Y(_0659_),
    .A(net444),
    .B(_0658_));
 sg13g2_o21ai_1 _2544_ (.B1(_0659_),
    .Y(_0262_),
    .A1(net444),
    .A2(\serialize.n433[1] ));
 sg13g2_nand4_1 _2545_ (.B(\videogen.fancy_shader.video_y[8] ),
    .C(\videogen.fancy_shader.video_y[7] ),
    .A(_0632_),
    .Y(_0660_),
    .D(\videogen.fancy_shader.video_y[6] ));
 sg13g2_nor2_1 _2546_ (.A(_0633_),
    .B(_0660_),
    .Y(_0661_));
 sg13g2_nand2b_1 _2547_ (.Y(_0662_),
    .B(_0661_),
    .A_N(\videogen.fancy_shader.video_y[4] ));
 sg13g2_nor2_1 _2548_ (.A(net608),
    .B(net609),
    .Y(_0663_));
 sg13g2_nor4_1 _2549_ (.A(\videogen.fancy_shader.video_y[3] ),
    .B(\videogen.fancy_shader.video_y[2] ),
    .C(net608),
    .D(net609),
    .Y(_0664_));
 sg13g2_nor2b_2 _2550_ (.A(_0662_),
    .B_N(_0664_),
    .Y(_0665_));
 sg13g2_nor2b_1 _2551_ (.A(\videogen.fancy_shader.video_x[8] ),
    .B_N(\videogen.fancy_shader.video_x[9] ),
    .Y(_0666_));
 sg13g2_and2_1 _2552_ (.A(net629),
    .B(_0666_),
    .X(_0667_));
 sg13g2_nor3_1 _2553_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(\videogen.fancy_shader.video_x[5] ),
    .C(\videogen.fancy_shader.video_x[4] ),
    .Y(_0668_));
 sg13g2_nor4_1 _2554_ (.A(\videogen.fancy_shader.video_x[3] ),
    .B(\videogen.fancy_shader.video_x[2] ),
    .C(\videogen.fancy_shader.video_x[1] ),
    .D(net630),
    .Y(_0669_));
 sg13g2_and3_2 _2555_ (.X(_0670_),
    .A(_0667_),
    .B(_0668_),
    .C(_0669_));
 sg13g2_nand3_1 _2556_ (.B(_0668_),
    .C(_0669_),
    .A(_0667_),
    .Y(_0671_));
 sg13g2_nor2_2 _2557_ (.A(_0665_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_nand2_2 _2558_ (.Y(_0673_),
    .A(net600),
    .B(_0672_));
 sg13g2_nor2_2 _2559_ (.A(net625),
    .B(net626),
    .Y(_0674_));
 sg13g2_or2_1 _2560_ (.X(_0675_),
    .B(net626),
    .A(net624));
 sg13g2_nor3_2 _2561_ (.A(net614),
    .B(net619),
    .C(net583),
    .Y(_0676_));
 sg13g2_a21oi_1 _2562_ (.A1(net592),
    .A2(_0674_),
    .Y(_0677_),
    .B1(net596));
 sg13g2_nor2_2 _2563_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_and2_1 _2564_ (.A(net543),
    .B(_0678_),
    .X(_0679_));
 sg13g2_nand2_2 _2565_ (.Y(_0680_),
    .A(net543),
    .B(_0678_));
 sg13g2_and2_1 _2566_ (.A(_0637_),
    .B(_0676_),
    .X(_0681_));
 sg13g2_xnor2_1 _2567_ (.Y(_0682_),
    .A(net612),
    .B(_0676_));
 sg13g2_and2_1 _2568_ (.A(_0636_),
    .B(_0681_),
    .X(_0683_));
 sg13g2_xnor2_1 _2569_ (.Y(_0684_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .B(_0681_));
 sg13g2_inv_1 _2570_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_a21oi_2 _2571_ (.B1(_0685_),
    .Y(_0686_),
    .A2(_0672_),
    .A1(net600));
 sg13g2_nand2_2 _2572_ (.Y(_0687_),
    .A(_0682_),
    .B(_0686_));
 sg13g2_nor2_2 _2573_ (.A(_0679_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_nand2b_2 _2574_ (.Y(_0689_),
    .B(_0680_),
    .A_N(_0687_));
 sg13g2_nand2_2 _2575_ (.Y(_0690_),
    .A(net624),
    .B(net626));
 sg13g2_and2_1 _2576_ (.A(net582),
    .B(net572),
    .X(_0691_));
 sg13g2_and2_1 _2577_ (.A(net543),
    .B(_0691_),
    .X(_0692_));
 sg13g2_nand2_1 _2578_ (.Y(_0693_),
    .A(net543),
    .B(_0691_));
 sg13g2_xnor2_1 _2579_ (.Y(_0694_),
    .A(net619),
    .B(_0674_));
 sg13g2_and2_1 _2580_ (.A(net543),
    .B(_0694_),
    .X(_0695_));
 sg13g2_nor2_1 _2581_ (.A(_0692_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_a21oi_2 _2582_ (.B1(_0649_),
    .Y(_0697_),
    .A2(net543),
    .A1(net626));
 sg13g2_and2_1 _2583_ (.A(_0696_),
    .B(_0697_),
    .X(_0698_));
 sg13g2_nand2_2 _2584_ (.Y(_0699_),
    .A(_0696_),
    .B(_0697_));
 sg13g2_nor2_2 _2585_ (.A(_0689_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_mux2_1 _2586_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .A1(net752),
    .S(_0700_),
    .X(_0631_));
 sg13g2_mux2_1 _2587_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .A1(net762),
    .S(_0700_),
    .X(_0630_));
 sg13g2_mux2_1 _2588_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .A1(net772),
    .S(_0700_),
    .X(_0629_));
 sg13g2_mux2_1 _2589_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .A1(net782),
    .S(_0700_),
    .X(_0628_));
 sg13g2_nand2_2 _2590_ (.Y(_0701_),
    .A(net600),
    .B(_0695_));
 sg13g2_nor2_2 _2591_ (.A(net588),
    .B(_0701_),
    .Y(_0702_));
 sg13g2_nand3_1 _2592_ (.B(_0674_),
    .C(_0695_),
    .A(\videogen.mem_read ),
    .Y(_0703_));
 sg13g2_nand2_2 _2593_ (.Y(_0704_),
    .A(_0688_),
    .B(_0702_));
 sg13g2_mux2_1 _2594_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .S(_0704_),
    .X(_0609_));
 sg13g2_mux2_1 _2595_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .S(_0704_),
    .X(_0608_));
 sg13g2_mux2_1 _2596_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ),
    .S(_0704_),
    .X(_0607_));
 sg13g2_mux2_1 _2597_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .S(_0704_),
    .X(_0606_));
 sg13g2_nand3_1 _2598_ (.B(_0682_),
    .C(_0685_),
    .A(net543),
    .Y(_0705_));
 sg13g2_nor2_2 _2599_ (.A(_0680_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_inv_1 _2600_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_nand2_2 _2601_ (.Y(_0708_),
    .A(_0698_),
    .B(_0706_));
 sg13g2_mux2_1 _2602_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .S(_0708_),
    .X(_0605_));
 sg13g2_mux2_1 _2603_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .S(_0708_),
    .X(_0604_));
 sg13g2_mux2_1 _2604_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .S(_0708_),
    .X(_0603_));
 sg13g2_mux2_1 _2605_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .S(_0708_),
    .X(_0602_));
 sg13g2_nand3_1 _2606_ (.B(net600),
    .C(net543),
    .A(net626),
    .Y(_0709_));
 sg13g2_nor3_2 _2607_ (.A(net619),
    .B(_0693_),
    .C(_0709_),
    .Y(_0710_));
 sg13g2_nand2_2 _2608_ (.Y(_0711_),
    .A(_0688_),
    .B(_0710_));
 sg13g2_mux2_1 _2609_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ),
    .S(_0711_),
    .X(_0601_));
 sg13g2_mux2_1 _2610_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .S(_0711_),
    .X(_0600_));
 sg13g2_mux2_1 _2611_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .S(_0711_),
    .X(_0599_));
 sg13g2_mux2_1 _2612_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ),
    .S(_0711_),
    .X(_0598_));
 sg13g2_nand2b_2 _2613_ (.Y(_0712_),
    .B(_0686_),
    .A_N(_0682_));
 sg13g2_nor2_2 _2614_ (.A(_0680_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_inv_1 _2615_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_and3_2 _2616_ (.X(_0715_),
    .A(net592),
    .B(_0692_),
    .C(_0697_));
 sg13g2_nand2_2 _2617_ (.Y(_0716_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_mux2_1 _2618_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .S(_0716_),
    .X(_0597_));
 sg13g2_mux2_1 _2619_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .S(_0716_),
    .X(_0596_));
 sg13g2_mux2_1 _2620_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .S(_0716_),
    .X(_0595_));
 sg13g2_mux2_1 _2621_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .S(_0716_),
    .X(_0594_));
 sg13g2_nor2_2 _2622_ (.A(net578),
    .B(_0701_),
    .Y(_0717_));
 sg13g2_or2_1 _2623_ (.X(_0718_),
    .B(_0701_),
    .A(net577));
 sg13g2_nand2_2 _2624_ (.Y(_0719_),
    .A(_0713_),
    .B(_0717_));
 sg13g2_mux2_1 _2625_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .S(_0719_),
    .X(_0593_));
 sg13g2_mux2_1 _2626_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .S(_0719_),
    .X(_0592_));
 sg13g2_mux2_1 _2627_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .S(_0719_),
    .X(_0591_));
 sg13g2_mux2_1 _2628_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .S(_0719_),
    .X(_0590_));
 sg13g2_nor2_2 _2629_ (.A(_0680_),
    .B(_0687_),
    .Y(_0720_));
 sg13g2_or2_1 _2630_ (.X(_0721_),
    .B(_0687_),
    .A(_0680_));
 sg13g2_and2_1 _2631_ (.A(_0715_),
    .B(_0720_),
    .X(_0722_));
 sg13g2_mux2_1 _2632_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .A1(net754),
    .S(_0722_),
    .X(_0589_));
 sg13g2_mux2_1 _2633_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .A1(net764),
    .S(_0722_),
    .X(_0588_));
 sg13g2_mux2_1 _2634_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .A1(net774),
    .S(_0722_),
    .X(_0587_));
 sg13g2_mux2_1 _2635_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .A1(net784),
    .S(_0722_),
    .X(_0586_));
 sg13g2_or3_1 _2636_ (.A(net592),
    .B(_0693_),
    .C(_0709_),
    .X(_0723_));
 sg13g2_nor2_2 _2637_ (.A(_0714_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_mux2_1 _2638_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .A1(net755),
    .S(_0724_),
    .X(_0585_));
 sg13g2_mux2_1 _2639_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .A1(net770),
    .S(_0724_),
    .X(_0584_));
 sg13g2_mux2_1 _2640_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .A1(net775),
    .S(_0724_),
    .X(_0583_));
 sg13g2_mux2_1 _2641_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .A1(net789),
    .S(_0724_),
    .X(_0582_));
 sg13g2_nand3_1 _2642_ (.B(_0692_),
    .C(_0697_),
    .A(net619),
    .Y(_0725_));
 sg13g2_nor2_2 _2643_ (.A(_0714_),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_mux2_1 _2644_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .A1(net755),
    .S(_0726_),
    .X(_0581_));
 sg13g2_mux2_1 _2645_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .A1(net770),
    .S(_0726_),
    .X(_0580_));
 sg13g2_mux2_1 _2646_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .A1(net775),
    .S(_0726_),
    .X(_0579_));
 sg13g2_mux2_1 _2647_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .A1(net789),
    .S(_0726_),
    .X(_0578_));
 sg13g2_nor3_2 _2648_ (.A(_0692_),
    .B(_0695_),
    .C(_0709_),
    .Y(_0727_));
 sg13g2_nand4_1 _2649_ (.B(net600),
    .C(_0673_),
    .A(net626),
    .Y(_0728_),
    .D(_0696_));
 sg13g2_nand2_2 _2650_ (.Y(_0729_),
    .A(_0713_),
    .B(_0727_));
 sg13g2_mux2_1 _2651_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .S(_0729_),
    .X(_0577_));
 sg13g2_mux2_1 _2652_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .S(_0729_),
    .X(_0576_));
 sg13g2_mux2_1 _2653_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .S(_0729_),
    .X(_0575_));
 sg13g2_mux2_1 _2654_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .S(_0729_),
    .X(_0574_));
 sg13g2_nand2_2 _2655_ (.Y(_0730_),
    .A(_0698_),
    .B(_0713_));
 sg13g2_mux2_1 _2656_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .S(_0730_),
    .X(_0573_));
 sg13g2_mux2_1 _2657_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .S(_0730_),
    .X(_0572_));
 sg13g2_mux2_1 _2658_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .S(_0730_),
    .X(_0571_));
 sg13g2_mux2_1 _2659_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .S(_0730_),
    .X(_0570_));
 sg13g2_nor2_2 _2660_ (.A(_0679_),
    .B(_0712_),
    .Y(_0731_));
 sg13g2_nand2_2 _2661_ (.Y(_0732_),
    .A(_0710_),
    .B(_0731_));
 sg13g2_mux2_1 _2662_ (.A0(net756),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .S(_0732_),
    .X(_0569_));
 sg13g2_mux2_1 _2663_ (.A0(net762),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .S(_0732_),
    .X(_0568_));
 sg13g2_mux2_1 _2664_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .S(_0732_),
    .X(_0567_));
 sg13g2_mux2_1 _2665_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ),
    .S(_0732_),
    .X(_0566_));
 sg13g2_nand2_2 _2666_ (.Y(_0733_),
    .A(_0715_),
    .B(_0731_));
 sg13g2_mux2_1 _2667_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .S(_0733_),
    .X(_0565_));
 sg13g2_mux2_1 _2668_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .S(_0733_),
    .X(_0564_));
 sg13g2_mux2_1 _2669_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .S(_0733_),
    .X(_0563_));
 sg13g2_mux2_1 _2670_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .S(_0733_),
    .X(_0562_));
 sg13g2_nand2_2 _2671_ (.Y(_0734_),
    .A(_0717_),
    .B(_0731_));
 sg13g2_mux2_1 _2672_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .S(_0734_),
    .X(_0561_));
 sg13g2_mux2_1 _2673_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .S(_0734_),
    .X(_0560_));
 sg13g2_mux2_1 _2674_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .S(_0734_),
    .X(_0559_));
 sg13g2_mux2_1 _2675_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ),
    .S(_0734_),
    .X(_0558_));
 sg13g2_nand2_2 _2676_ (.Y(_0735_),
    .A(_0702_),
    .B(_0731_));
 sg13g2_mux2_1 _2677_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ),
    .S(_0735_),
    .X(_0557_));
 sg13g2_mux2_1 _2678_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .S(_0735_),
    .X(_0556_));
 sg13g2_mux2_1 _2679_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ),
    .S(_0735_),
    .X(_0555_));
 sg13g2_mux2_1 _2680_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .S(_0735_),
    .X(_0554_));
 sg13g2_nor2b_2 _2681_ (.A(_0723_),
    .B_N(_0731_),
    .Y(_0736_));
 sg13g2_mux2_1 _2682_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .A1(net755),
    .S(_0736_),
    .X(_0553_));
 sg13g2_mux2_1 _2683_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .A1(net766),
    .S(_0736_),
    .X(_0552_));
 sg13g2_mux2_1 _2684_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .A1(net775),
    .S(_0736_),
    .X(_0551_));
 sg13g2_mux2_1 _2685_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .A1(net786),
    .S(_0736_),
    .X(_0550_));
 sg13g2_nand2_2 _2686_ (.Y(_0737_),
    .A(_0717_),
    .B(_0720_));
 sg13g2_mux2_1 _2687_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .S(_0737_),
    .X(_0549_));
 sg13g2_mux2_1 _2688_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .S(_0737_),
    .X(_0548_));
 sg13g2_mux2_1 _2689_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .S(_0737_),
    .X(_0547_));
 sg13g2_mux2_1 _2690_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .S(_0737_),
    .X(_0546_));
 sg13g2_nand2_2 _2691_ (.Y(_0738_),
    .A(_0727_),
    .B(_0731_));
 sg13g2_mux2_1 _2692_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .S(_0738_),
    .X(_0545_));
 sg13g2_mux2_1 _2693_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .S(_0738_),
    .X(_0544_));
 sg13g2_mux2_1 _2694_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .S(_0738_),
    .X(_0543_));
 sg13g2_mux2_1 _2695_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ),
    .S(_0738_),
    .X(_0542_));
 sg13g2_nand2_2 _2696_ (.Y(_0739_),
    .A(_0698_),
    .B(_0731_));
 sg13g2_mux2_1 _2697_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .S(_0739_),
    .X(_0541_));
 sg13g2_mux2_1 _2698_ (.A0(net766),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .S(_0739_),
    .X(_0540_));
 sg13g2_mux2_1 _2699_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .S(_0739_),
    .X(_0539_));
 sg13g2_mux2_1 _2700_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ),
    .S(_0739_),
    .X(_0538_));
 sg13g2_nand2_2 _2701_ (.Y(_0740_),
    .A(_0706_),
    .B(_0710_));
 sg13g2_mux2_1 _2702_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .S(_0740_),
    .X(_0537_));
 sg13g2_mux2_1 _2703_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .S(_0740_),
    .X(_0536_));
 sg13g2_mux2_1 _2704_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .S(_0740_),
    .X(_0535_));
 sg13g2_mux2_1 _2705_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .S(_0740_),
    .X(_0534_));
 sg13g2_nand2_2 _2706_ (.Y(_0741_),
    .A(_0706_),
    .B(_0715_));
 sg13g2_mux2_1 _2707_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .S(_0741_),
    .X(_0533_));
 sg13g2_mux2_1 _2708_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .S(_0741_),
    .X(_0532_));
 sg13g2_mux2_1 _2709_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .S(_0741_),
    .X(_0531_));
 sg13g2_mux2_1 _2710_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .S(_0741_),
    .X(_0530_));
 sg13g2_nand2_2 _2711_ (.Y(_0742_),
    .A(_0706_),
    .B(_0717_));
 sg13g2_mux2_1 _2712_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .S(_0742_),
    .X(_0529_));
 sg13g2_mux2_1 _2713_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .S(_0742_),
    .X(_0528_));
 sg13g2_mux2_1 _2714_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .S(_0742_),
    .X(_0527_));
 sg13g2_mux2_1 _2715_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .S(_0742_),
    .X(_0526_));
 sg13g2_nand2_2 _2716_ (.Y(_0743_),
    .A(_0702_),
    .B(_0706_));
 sg13g2_mux2_1 _2717_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .S(_0743_),
    .X(_0525_));
 sg13g2_mux2_1 _2718_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .S(_0743_),
    .X(_0524_));
 sg13g2_mux2_1 _2719_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ),
    .S(_0743_),
    .X(_0523_));
 sg13g2_mux2_1 _2720_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ),
    .S(_0743_),
    .X(_0522_));
 sg13g2_nor2_2 _2721_ (.A(_0707_),
    .B(_0723_),
    .Y(_0744_));
 sg13g2_mux2_1 _2722_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .A1(net759),
    .S(_0744_),
    .X(_0521_));
 sg13g2_mux2_1 _2723_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .A1(net769),
    .S(_0744_),
    .X(_0520_));
 sg13g2_mux2_1 _2724_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .A1(net780),
    .S(_0744_),
    .X(_0519_));
 sg13g2_mux2_1 _2725_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .A1(net790),
    .S(_0744_),
    .X(_0518_));
 sg13g2_nor2_2 _2726_ (.A(_0707_),
    .B(_0725_),
    .Y(_0745_));
 sg13g2_mux2_1 _2727_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .A1(net759),
    .S(_0745_),
    .X(_0517_));
 sg13g2_mux2_1 _2728_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .A1(net769),
    .S(_0745_),
    .X(_0516_));
 sg13g2_mux2_1 _2729_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .A1(net780),
    .S(_0745_),
    .X(_0515_));
 sg13g2_mux2_1 _2730_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .A1(net790),
    .S(_0745_),
    .X(_0514_));
 sg13g2_nand2_2 _2731_ (.Y(_0746_),
    .A(_0706_),
    .B(_0727_));
 sg13g2_mux2_1 _2732_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .S(_0746_),
    .X(_0513_));
 sg13g2_mux2_1 _2733_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .S(_0746_),
    .X(_0512_));
 sg13g2_mux2_1 _2734_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .S(_0746_),
    .X(_0511_));
 sg13g2_mux2_1 _2735_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .S(_0746_),
    .X(_0510_));
 sg13g2_nand2_2 _2736_ (.Y(_0747_),
    .A(_0702_),
    .B(_0720_));
 sg13g2_mux2_1 _2737_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ),
    .S(_0747_),
    .X(_0509_));
 sg13g2_mux2_1 _2738_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .S(_0747_),
    .X(_0508_));
 sg13g2_mux2_1 _2739_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .S(_0747_),
    .X(_0507_));
 sg13g2_mux2_1 _2740_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .S(_0747_),
    .X(_0506_));
 sg13g2_nand2_2 _2741_ (.Y(_0748_),
    .A(_0688_),
    .B(_0727_));
 sg13g2_mux2_1 _2742_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .S(_0748_),
    .X(_0496_));
 sg13g2_mux2_1 _2743_ (.A0(net762),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .S(_0748_),
    .X(_0495_));
 sg13g2_mux2_1 _2744_ (.A0(net772),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .S(_0748_),
    .X(_0494_));
 sg13g2_mux2_1 _2745_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .S(_0748_),
    .X(_0493_));
 sg13g2_nor2_2 _2746_ (.A(_0689_),
    .B(_0723_),
    .Y(_0749_));
 sg13g2_mux2_1 _2747_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .A1(net752),
    .S(_0749_),
    .X(_0492_));
 sg13g2_mux2_1 _2748_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .A1(net762),
    .S(_0749_),
    .X(_0491_));
 sg13g2_mux2_1 _2749_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .A1(net772),
    .S(_0749_),
    .X(_0490_));
 sg13g2_mux2_1 _2750_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .A1(net782),
    .S(_0749_),
    .X(_0489_));
 sg13g2_nand2_2 _2751_ (.Y(_0750_),
    .A(_0710_),
    .B(_0713_));
 sg13g2_mux2_1 _2752_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ),
    .S(_0750_),
    .X(_0488_));
 sg13g2_mux2_1 _2753_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .S(_0750_),
    .X(_0487_));
 sg13g2_mux2_1 _2754_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ),
    .S(_0750_),
    .X(_0486_));
 sg13g2_mux2_1 _2755_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ),
    .S(_0750_),
    .X(_0485_));
 sg13g2_nor2_2 _2756_ (.A(_0679_),
    .B(_0705_),
    .Y(_0751_));
 sg13g2_nand2_2 _2757_ (.Y(_0752_),
    .A(_0715_),
    .B(_0751_));
 sg13g2_mux2_1 _2758_ (.A0(net756),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .S(_0752_),
    .X(_0484_));
 sg13g2_mux2_1 _2759_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .S(_0752_),
    .X(_0483_));
 sg13g2_mux2_1 _2760_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ),
    .S(_0752_),
    .X(_0482_));
 sg13g2_mux2_1 _2761_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ),
    .S(_0752_),
    .X(_0481_));
 sg13g2_nand2_2 _2762_ (.Y(_0753_),
    .A(_0710_),
    .B(_0751_));
 sg13g2_mux2_1 _2763_ (.A0(net756),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .S(_0753_),
    .X(_0480_));
 sg13g2_mux2_1 _2764_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .S(_0753_),
    .X(_0479_));
 sg13g2_mux2_1 _2765_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .S(_0753_),
    .X(_0478_));
 sg13g2_mux2_1 _2766_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .S(_0753_),
    .X(_0477_));
 sg13g2_nand2_2 _2767_ (.Y(_0754_),
    .A(_0710_),
    .B(_0720_));
 sg13g2_mux2_1 _2768_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .S(_0754_),
    .X(_0476_));
 sg13g2_mux2_1 _2769_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .S(_0754_),
    .X(_0475_));
 sg13g2_mux2_1 _2770_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ),
    .S(_0754_),
    .X(_0474_));
 sg13g2_mux2_1 _2771_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ),
    .S(_0754_),
    .X(_0473_));
 sg13g2_nand2_2 _2772_ (.Y(_0755_),
    .A(_0717_),
    .B(_0751_));
 sg13g2_mux2_1 _2773_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .S(_0755_),
    .X(_0472_));
 sg13g2_mux2_1 _2774_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .S(_0755_),
    .X(_0471_));
 sg13g2_mux2_1 _2775_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .S(_0755_),
    .X(_0470_));
 sg13g2_mux2_1 _2776_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .S(_0755_),
    .X(_0469_));
 sg13g2_nand2_2 _2777_ (.Y(_0756_),
    .A(_0702_),
    .B(_0751_));
 sg13g2_mux2_1 _2778_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .S(_0756_),
    .X(_0468_));
 sg13g2_mux2_1 _2779_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .S(_0756_),
    .X(_0467_));
 sg13g2_mux2_1 _2780_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .S(_0756_),
    .X(_0466_));
 sg13g2_mux2_1 _2781_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .S(_0756_),
    .X(_0465_));
 sg13g2_nor2b_2 _2782_ (.A(_0723_),
    .B_N(_0751_),
    .Y(_0757_));
 sg13g2_mux2_1 _2783_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ),
    .A1(net756),
    .S(_0757_),
    .X(_0464_));
 sg13g2_mux2_1 _2784_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .A1(net771),
    .S(_0757_),
    .X(_0463_));
 sg13g2_mux2_1 _2785_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .A1(net778),
    .S(_0757_),
    .X(_0462_));
 sg13g2_mux2_1 _2786_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .A1(net788),
    .S(_0757_),
    .X(_0461_));
 sg13g2_nor2b_2 _2787_ (.A(_0725_),
    .B_N(_0751_),
    .Y(_0758_));
 sg13g2_mux2_1 _2788_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .A1(net757),
    .S(_0758_),
    .X(_0460_));
 sg13g2_mux2_1 _2789_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .A1(net767),
    .S(_0758_),
    .X(_0459_));
 sg13g2_mux2_1 _2790_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .A1(net778),
    .S(_0758_),
    .X(_0458_));
 sg13g2_mux2_1 _2791_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ),
    .A1(net788),
    .S(_0758_),
    .X(_0457_));
 sg13g2_nand2_2 _2792_ (.Y(_0759_),
    .A(_0727_),
    .B(_0751_));
 sg13g2_mux2_1 _2793_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .S(_0759_),
    .X(_0456_));
 sg13g2_mux2_1 _2794_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .S(_0759_),
    .X(_0455_));
 sg13g2_mux2_1 _2795_ (.A0(net778),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .S(_0759_),
    .X(_0454_));
 sg13g2_mux2_1 _2796_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ),
    .S(_0759_),
    .X(_0453_));
 sg13g2_nand2_2 _2797_ (.Y(_0760_),
    .A(_0698_),
    .B(_0751_));
 sg13g2_mux2_1 _2798_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ),
    .S(_0760_),
    .X(_0452_));
 sg13g2_mux2_1 _2799_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .S(_0760_),
    .X(_0451_));
 sg13g2_mux2_1 _2800_ (.A0(net778),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .S(_0760_),
    .X(_0450_));
 sg13g2_mux2_1 _2801_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .S(_0760_),
    .X(_0449_));
 sg13g2_o21ai_1 _2802_ (.B1(_0673_),
    .Y(_0761_),
    .A1(_0682_),
    .A2(_0684_));
 sg13g2_nand2_2 _2803_ (.Y(_0762_),
    .A(_0679_),
    .B(_0761_));
 sg13g2_inv_1 _2804_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_nand2_2 _2805_ (.Y(_0764_),
    .A(_0710_),
    .B(_0763_));
 sg13g2_mux2_1 _2806_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .S(_0764_),
    .X(_0448_));
 sg13g2_mux2_1 _2807_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .S(_0764_),
    .X(_0447_));
 sg13g2_mux2_1 _2808_ (.A0(net778),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .S(_0764_),
    .X(_0446_));
 sg13g2_mux2_1 _2809_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .S(_0764_),
    .X(_0445_));
 sg13g2_nor2_2 _2810_ (.A(_0721_),
    .B(_0723_),
    .Y(_0765_));
 sg13g2_mux2_1 _2811_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .A1(net753),
    .S(_0765_),
    .X(_0444_));
 sg13g2_mux2_1 _2812_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .A1(net764),
    .S(_0765_),
    .X(_0443_));
 sg13g2_mux2_1 _2813_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .A1(net773),
    .S(_0765_),
    .X(_0442_));
 sg13g2_mux2_1 _2814_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .A1(net785),
    .S(_0765_),
    .X(_0441_));
 sg13g2_nor2_2 _2815_ (.A(_0718_),
    .B(_0762_),
    .Y(_0766_));
 sg13g2_mux2_1 _2816_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .A1(net757),
    .S(_0766_),
    .X(_0440_));
 sg13g2_mux2_1 _2817_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .A1(net767),
    .S(_0766_),
    .X(_0439_));
 sg13g2_mux2_1 _2818_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .A1(net778),
    .S(_0766_),
    .X(_0438_));
 sg13g2_mux2_1 _2819_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .A1(net788),
    .S(_0766_),
    .X(_0437_));
 sg13g2_nor2_2 _2820_ (.A(_0703_),
    .B(_0762_),
    .Y(_0767_));
 sg13g2_mux2_1 _2821_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .A1(net757),
    .S(_0767_),
    .X(_0436_));
 sg13g2_mux2_1 _2822_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .A1(net767),
    .S(_0767_),
    .X(_0435_));
 sg13g2_mux2_1 _2823_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ),
    .A1(net778),
    .S(_0767_),
    .X(_0434_));
 sg13g2_mux2_1 _2824_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .A1(net788),
    .S(_0767_),
    .X(_0433_));
 sg13g2_nor2_2 _2825_ (.A(_0723_),
    .B(_0762_),
    .Y(_0768_));
 sg13g2_mux2_1 _2826_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .A1(net753),
    .S(_0768_),
    .X(_0432_));
 sg13g2_mux2_1 _2827_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .A1(net768),
    .S(_0768_),
    .X(_0431_));
 sg13g2_mux2_1 _2828_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .A1(net773),
    .S(_0768_),
    .X(_0430_));
 sg13g2_mux2_1 _2829_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ),
    .A1(net783),
    .S(_0768_),
    .X(_0429_));
 sg13g2_nor2_2 _2830_ (.A(_0725_),
    .B(_0762_),
    .Y(_0769_));
 sg13g2_mux2_1 _2831_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .A1(net753),
    .S(_0769_),
    .X(_0428_));
 sg13g2_mux2_1 _2832_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .A1(net763),
    .S(_0769_),
    .X(_0427_));
 sg13g2_mux2_1 _2833_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .A1(net773),
    .S(_0769_),
    .X(_0426_));
 sg13g2_mux2_1 _2834_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .A1(net783),
    .S(_0769_),
    .X(_0425_));
 sg13g2_nor2_2 _2835_ (.A(_0728_),
    .B(_0762_),
    .Y(_0770_));
 sg13g2_mux2_1 _2836_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .A1(net753),
    .S(_0770_),
    .X(_0424_));
 sg13g2_mux2_1 _2837_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .A1(net763),
    .S(_0770_),
    .X(_0423_));
 sg13g2_mux2_1 _2838_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .A1(net773),
    .S(_0770_),
    .X(_0422_));
 sg13g2_mux2_1 _2839_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .A1(net783),
    .S(_0770_),
    .X(_0421_));
 sg13g2_nor2_2 _2840_ (.A(_0699_),
    .B(_0762_),
    .Y(_0771_));
 sg13g2_mux2_1 _2841_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .A1(net753),
    .S(_0771_),
    .X(_0420_));
 sg13g2_mux2_1 _2842_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .A1(net768),
    .S(_0771_),
    .X(_0419_));
 sg13g2_mux2_1 _2843_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .A1(net773),
    .S(_0771_),
    .X(_0418_));
 sg13g2_mux2_1 _2844_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ),
    .A1(net783),
    .S(_0771_),
    .X(_0417_));
 sg13g2_nand2_2 _2845_ (.Y(_0772_),
    .A(_0680_),
    .B(_0761_));
 sg13g2_inv_1 _2846_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_nand2_2 _2847_ (.Y(_0774_),
    .A(_0710_),
    .B(_0773_));
 sg13g2_mux2_1 _2848_ (.A0(net756),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .S(_0774_),
    .X(_0416_));
 sg13g2_mux2_1 _2849_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .S(_0774_),
    .X(_0415_));
 sg13g2_mux2_1 _2850_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .S(_0774_),
    .X(_0414_));
 sg13g2_mux2_1 _2851_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ),
    .S(_0774_),
    .X(_0413_));
 sg13g2_nand2_2 _2852_ (.Y(_0775_),
    .A(_0715_),
    .B(_0773_));
 sg13g2_mux2_1 _2853_ (.A0(net756),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .S(_0775_),
    .X(_0412_));
 sg13g2_mux2_1 _2854_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .S(_0775_),
    .X(_0411_));
 sg13g2_mux2_1 _2855_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ),
    .S(_0775_),
    .X(_0410_));
 sg13g2_mux2_1 _2856_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .S(_0775_),
    .X(_0409_));
 sg13g2_nor2_2 _2857_ (.A(_0718_),
    .B(_0772_),
    .Y(_0776_));
 sg13g2_mux2_1 _2858_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .A1(net756),
    .S(_0776_),
    .X(_0408_));
 sg13g2_mux2_1 _2859_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .A1(net768),
    .S(_0776_),
    .X(_0407_));
 sg13g2_mux2_1 _2860_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .A1(net777),
    .S(_0776_),
    .X(_0406_));
 sg13g2_mux2_1 _2861_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .A1(net787),
    .S(_0776_),
    .X(_0405_));
 sg13g2_nor2_2 _2862_ (.A(_0721_),
    .B(_0725_),
    .Y(_0777_));
 sg13g2_mux2_1 _2863_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .A1(net761),
    .S(_0777_),
    .X(_0404_));
 sg13g2_mux2_1 _2864_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .A1(net764),
    .S(_0777_),
    .X(_0403_));
 sg13g2_mux2_1 _2865_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .A1(net773),
    .S(_0777_),
    .X(_0402_));
 sg13g2_mux2_1 _2866_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .A1(net785),
    .S(_0777_),
    .X(_0401_));
 sg13g2_nor2_2 _2867_ (.A(_0723_),
    .B(_0772_),
    .Y(_0778_));
 sg13g2_mux2_1 _2868_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .A1(net752),
    .S(_0778_),
    .X(_0400_));
 sg13g2_mux2_1 _2869_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ),
    .A1(net762),
    .S(_0778_),
    .X(_0399_));
 sg13g2_mux2_1 _2870_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ),
    .A1(net772),
    .S(_0778_),
    .X(_0398_));
 sg13g2_mux2_1 _2871_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ),
    .A1(net782),
    .S(_0778_),
    .X(_0397_));
 sg13g2_nor2_2 _2872_ (.A(_0725_),
    .B(_0772_),
    .Y(_0779_));
 sg13g2_mux2_1 _2873_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .A1(net752),
    .S(_0779_),
    .X(_0396_));
 sg13g2_mux2_1 _2874_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .A1(net762),
    .S(_0779_),
    .X(_0395_));
 sg13g2_mux2_1 _2875_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .A1(net772),
    .S(_0779_),
    .X(_0394_));
 sg13g2_mux2_1 _2876_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .A1(net782),
    .S(_0779_),
    .X(_0393_));
 sg13g2_nor2_2 _2877_ (.A(_0728_),
    .B(_0772_),
    .Y(_0780_));
 sg13g2_mux2_1 _2878_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .A1(net752),
    .S(_0780_),
    .X(_0392_));
 sg13g2_mux2_1 _2879_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .A1(net762),
    .S(_0780_),
    .X(_0391_));
 sg13g2_mux2_1 _2880_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .A1(net772),
    .S(_0780_),
    .X(_0390_));
 sg13g2_mux2_1 _2881_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .A1(net783),
    .S(_0780_),
    .X(_0389_));
 sg13g2_nor2_2 _2882_ (.A(_0689_),
    .B(_0725_),
    .Y(_0781_));
 sg13g2_mux2_1 _2883_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .A1(net752),
    .S(_0781_),
    .X(_0345_));
 sg13g2_mux2_1 _2884_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .A1(net762),
    .S(_0781_),
    .X(_0344_));
 sg13g2_mux2_1 _2885_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .A1(net772),
    .S(_0781_),
    .X(_0343_));
 sg13g2_mux2_1 _2886_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .A1(net782),
    .S(_0781_),
    .X(_0342_));
 sg13g2_nand2_2 _2887_ (.Y(_0782_),
    .A(_0702_),
    .B(_0713_));
 sg13g2_mux2_1 _2888_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .S(_0782_),
    .X(_0341_));
 sg13g2_mux2_1 _2889_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .S(_0782_),
    .X(_0340_));
 sg13g2_mux2_1 _2890_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .S(_0782_),
    .X(_0339_));
 sg13g2_mux2_1 _2891_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .S(_0782_),
    .X(_0338_));
 sg13g2_nor2b_2 _2892_ (.A(_0725_),
    .B_N(_0731_),
    .Y(_0783_));
 sg13g2_mux2_1 _2893_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .A1(net755),
    .S(_0783_),
    .X(_0316_));
 sg13g2_mux2_1 _2894_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .A1(net766),
    .S(_0783_),
    .X(_0315_));
 sg13g2_mux2_1 _2895_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .A1(net776),
    .S(_0783_),
    .X(_0314_));
 sg13g2_mux2_1 _2896_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .A1(net786),
    .S(_0783_),
    .X(_0313_));
 sg13g2_nand2_2 _2897_ (.Y(_0784_),
    .A(_0688_),
    .B(_0717_));
 sg13g2_mux2_1 _2898_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .S(_0784_),
    .X(_0302_));
 sg13g2_mux2_1 _2899_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .S(_0784_),
    .X(_0301_));
 sg13g2_mux2_1 _2900_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .S(_0784_),
    .X(_0300_));
 sg13g2_mux2_1 _2901_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .S(_0784_),
    .X(_0299_));
 sg13g2_nand2_2 _2902_ (.Y(_0785_),
    .A(_0720_),
    .B(_0727_));
 sg13g2_mux2_1 _2903_ (.A0(net753),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .S(_0785_),
    .X(_0298_));
 sg13g2_mux2_1 _2904_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .S(_0785_),
    .X(_0297_));
 sg13g2_mux2_1 _2905_ (.A0(net773),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .S(_0785_),
    .X(_0296_));
 sg13g2_mux2_1 _2906_ (.A0(net785),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .S(_0785_),
    .X(_0295_));
 sg13g2_nand2_2 _2907_ (.Y(_0786_),
    .A(_0688_),
    .B(_0715_));
 sg13g2_mux2_1 _2908_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .S(_0786_),
    .X(_0294_));
 sg13g2_mux2_1 _2909_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .S(_0786_),
    .X(_0293_));
 sg13g2_mux2_1 _2910_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .S(_0786_),
    .X(_0292_));
 sg13g2_mux2_1 _2911_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .S(_0786_),
    .X(_0291_));
 sg13g2_nor2_2 _2912_ (.A(_0703_),
    .B(_0772_),
    .Y(_0787_));
 sg13g2_mux2_1 _2913_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .A1(net756),
    .S(_0787_),
    .X(_0290_));
 sg13g2_mux2_1 _2914_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .A1(net768),
    .S(_0787_),
    .X(_0289_));
 sg13g2_mux2_1 _2915_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .A1(net777),
    .S(_0787_),
    .X(_0288_));
 sg13g2_mux2_1 _2916_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .A1(net787),
    .S(_0787_),
    .X(_0287_));
 sg13g2_nor2_2 _2917_ (.A(_0699_),
    .B(_0721_),
    .Y(_0788_));
 sg13g2_mux2_1 _2918_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .A1(net753),
    .S(_0788_),
    .X(_0286_));
 sg13g2_mux2_1 _2919_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .A1(net763),
    .S(_0788_),
    .X(_0285_));
 sg13g2_mux2_1 _2920_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .A1(net776),
    .S(_0788_),
    .X(_0284_));
 sg13g2_mux2_1 _2921_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .A1(net785),
    .S(_0788_),
    .X(_0283_));
 sg13g2_nor2_2 _2922_ (.A(_0699_),
    .B(_0772_),
    .Y(_0789_));
 sg13g2_mux2_1 _2923_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ),
    .A1(net752),
    .S(_0789_),
    .X(_0282_));
 sg13g2_mux2_1 _2924_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .A1(net763),
    .S(_0789_),
    .X(_0281_));
 sg13g2_mux2_1 _2925_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ),
    .A1(net772),
    .S(_0789_),
    .X(_0280_));
 sg13g2_mux2_1 _2926_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .A1(net783),
    .S(_0789_),
    .X(_0279_));
 sg13g2_nand2_2 _2927_ (.Y(_0790_),
    .A(_0715_),
    .B(_0763_));
 sg13g2_mux2_1 _2928_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .S(_0790_),
    .X(_0270_));
 sg13g2_mux2_1 _2929_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .S(_0790_),
    .X(_0269_));
 sg13g2_mux2_1 _2930_ (.A0(net778),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .S(_0790_),
    .X(_0268_));
 sg13g2_mux2_1 _2931_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ),
    .S(_0790_),
    .X(_0267_));
 sg13g2_and2_1 _2932_ (.A(\videogen.fancy_shader.video_x[8] ),
    .B(\videogen.fancy_shader.video_x[9] ),
    .X(_0791_));
 sg13g2_nor4_2 _2933_ (.A(\videogen.fancy_shader.video_y[9] ),
    .B(_0661_),
    .C(_0667_),
    .Y(_0792_),
    .D(_0791_));
 sg13g2_and2_1 _2934_ (.A(net793),
    .B(_0792_),
    .X(_0371_));
 sg13g2_nand2b_2 _2935_ (.Y(_0793_),
    .B(net793),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ));
 sg13g2_inv_2 _2936_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_and3_2 _2937_ (.X(_0795_),
    .A(\videogen.fancy_shader.video_x[2] ),
    .B(\videogen.fancy_shader.video_x[1] ),
    .C(net630));
 sg13g2_and2_1 _2938_ (.A(\videogen.fancy_shader.video_x[3] ),
    .B(_0795_),
    .X(_0796_));
 sg13g2_nand2_1 _2939_ (.Y(_0797_),
    .A(\videogen.fancy_shader.video_x[3] ),
    .B(_0795_));
 sg13g2_and2_1 _2940_ (.A(\videogen.fancy_shader.video_x[4] ),
    .B(_0796_),
    .X(_0798_));
 sg13g2_and2_1 _2941_ (.A(\videogen.fancy_shader.video_x[5] ),
    .B(_0798_),
    .X(_0799_));
 sg13g2_and2_1 _2942_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(_0799_),
    .X(_0800_));
 sg13g2_nor2b_1 _2943_ (.A(net629),
    .B_N(_0666_),
    .Y(_0801_));
 sg13g2_and2_1 _2944_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .B(_0792_),
    .X(_0802_));
 sg13g2_nand2_1 _2945_ (.Y(_0803_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ));
 sg13g2_nor3_2 _2946_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_nor2_1 _2947_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .Y(_0805_));
 sg13g2_and3_1 _2948_ (.X(_0806_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .B(_0804_),
    .C(_0805_));
 sg13g2_a22oi_1 _2949_ (.Y(_0807_),
    .B1(_0802_),
    .B2(_0806_),
    .A2(_0801_),
    .A1(_0800_));
 sg13g2_nand2b_1 _2950_ (.Y(_0808_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ),
    .A_N(_0792_));
 sg13g2_or2_1 _2951_ (.X(_0809_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.state[3] ),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ));
 sg13g2_nand2_1 _2952_ (.Y(_0810_),
    .A(net793),
    .B(_0809_));
 sg13g2_nand4_1 _2953_ (.B(_0807_),
    .C(_0808_),
    .A(net793),
    .Y(_0811_),
    .D(_0809_));
 sg13g2_a21oi_1 _2954_ (.A1(_0794_),
    .A2(_0811_),
    .Y(_0002_),
    .B1(_0371_));
 sg13g2_o21ai_1 _2955_ (.B1(_0792_),
    .Y(_0812_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ),
    .A2(_0807_));
 sg13g2_a21oi_1 _2956_ (.A1(_0649_),
    .A2(_0812_),
    .Y(_0003_),
    .B1(net747));
 sg13g2_nor3_2 _2957_ (.A(net429),
    .B(net413),
    .C(net446),
    .Y(\serialize.n410 ));
 sg13g2_a21o_2 _2958_ (.A2(_0804_),
    .A1(_0792_),
    .B1(\videogen.mem_read ),
    .X(\videogen.mem_row ));
 sg13g2_a21oi_2 _2959_ (.B1(_0649_),
    .Y(net8),
    .A2(_0671_),
    .A1(net627));
 sg13g2_a21oi_2 _2960_ (.B1(_0649_),
    .Y(net9),
    .A2(_0691_),
    .A1(_0671_));
 sg13g2_a21oi_2 _2961_ (.B1(_0649_),
    .Y(net10),
    .A2(_0694_),
    .A1(_0671_));
 sg13g2_a21oi_2 _2962_ (.B1(_0649_),
    .Y(net13),
    .A2(_0678_),
    .A1(_0671_));
 sg13g2_a21oi_2 _2963_ (.B1(_0649_),
    .Y(net14),
    .A2(_0682_),
    .A1(_0671_));
 sg13g2_a21oi_2 _2964_ (.B1(_0649_),
    .Y(net15),
    .A2(_0684_),
    .A1(_0671_));
 sg13g2_and2_1 _2965_ (.A(_0671_),
    .B(_0683_),
    .X(_0813_));
 sg13g2_and2_1 _2966_ (.A(net608),
    .B(net609),
    .X(_0814_));
 sg13g2_nand2_1 _2967_ (.Y(_0815_),
    .A(net608),
    .B(net609));
 sg13g2_nand3_1 _2968_ (.B(\videogen.fancy_shader.video_y[3] ),
    .C(\videogen.fancy_shader.video_y[2] ),
    .A(\videogen.fancy_shader.video_y[4] ),
    .Y(_0816_));
 sg13g2_nor4_1 _2969_ (.A(\videogen.fancy_shader.video_y[5] ),
    .B(_0660_),
    .C(_0815_),
    .D(_0816_),
    .Y(_0817_));
 sg13g2_nor2_2 _2970_ (.A(_0665_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_inv_1 _2971_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_o21ai_1 _2972_ (.B1(net600),
    .Y(_0820_),
    .A1(_0813_),
    .A2(_0818_));
 sg13g2_nor2_2 _2973_ (.A(_0670_),
    .B(_0683_),
    .Y(_0821_));
 sg13g2_and2_1 _2974_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0821_),
    .X(_0822_));
 sg13g2_xnor2_1 _2975_ (.Y(_0823_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0821_));
 sg13g2_a21oi_1 _2976_ (.A1(_0818_),
    .A2(_0823_),
    .Y(net16),
    .B1(_0820_));
 sg13g2_xnor2_1 _2977_ (.Y(_0824_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .B(_0822_));
 sg13g2_a21oi_1 _2978_ (.A1(_0818_),
    .A2(_0824_),
    .Y(net17),
    .B1(_0820_));
 sg13g2_and3_2 _2979_ (.X(_0825_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .C(_0822_));
 sg13g2_a21oi_1 _2980_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .A2(_0822_),
    .Y(_0826_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ));
 sg13g2_o21ai_1 _2981_ (.B1(_0818_),
    .Y(_0827_),
    .A1(_0825_),
    .A2(_0826_));
 sg13g2_nor2b_1 _2982_ (.A(_0820_),
    .B_N(_0827_),
    .Y(net18));
 sg13g2_xnor2_1 _2983_ (.Y(_0828_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B(_0825_));
 sg13g2_a21oi_1 _2984_ (.A1(_0818_),
    .A2(_0828_),
    .Y(net19),
    .B1(_0820_));
 sg13g2_nand3_1 _2985_ (.B(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .C(_0825_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .Y(_0829_));
 sg13g2_a21o_1 _2986_ (.A2(_0825_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .X(_0830_));
 sg13g2_a21oi_1 _2987_ (.A1(_0829_),
    .A2(_0830_),
    .Y(_0831_),
    .B1(_0819_));
 sg13g2_nor2_1 _2988_ (.A(_0820_),
    .B(_0831_),
    .Y(net20));
 sg13g2_or2_1 _2989_ (.X(_0832_),
    .B(_0829_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ));
 sg13g2_a21oi_1 _2990_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0829_),
    .Y(_0833_),
    .B1(_0819_));
 sg13g2_a21oi_1 _2991_ (.A1(_0832_),
    .A2(_0833_),
    .Y(net7),
    .B1(_0820_));
 sg13g2_mux2_1 _2992_ (.A0(\serialize.n461 ),
    .A1(\serialize.n459 ),
    .S(clknet_1_0__leaf_clk),
    .X(net4));
 sg13g2_mux2_1 _2993_ (.A0(\serialize.n458 ),
    .A1(\serialize.n456 ),
    .S(clknet_1_0__leaf_clk),
    .X(net3));
 sg13g2_mux2_1 _2994_ (.A0(\serialize.n455 ),
    .A1(\serialize.n453 ),
    .S(clknet_1_1__leaf_clk),
    .X(net5));
 sg13g2_mux2_1 _2995_ (.A0(\serialize.n452 ),
    .A1(\serialize.n450 ),
    .S(clknet_1_1__leaf_clk),
    .X(net6));
 sg13g2_nor2_1 _2996_ (.A(net413),
    .B(net695),
    .Y(\serialize.n433[0] ));
 sg13g2_nor2b_1 _2997_ (.A(net699),
    .B_N(net409),
    .Y(\serialize.n431[0] ));
 sg13g2_nor2b_1 _2998_ (.A(net699),
    .B_N(net408),
    .Y(\serialize.n431[1] ));
 sg13g2_nor2b_1 _2999_ (.A(net700),
    .B_N(net410),
    .Y(\serialize.n431[2] ));
 sg13g2_nor2b_1 _3000_ (.A(net700),
    .B_N(net411),
    .Y(\serialize.n431[3] ));
 sg13g2_nor2b_1 _3001_ (.A(net699),
    .B_N(net412),
    .Y(\serialize.n431[4] ));
 sg13g2_or2_1 _3002_ (.X(\serialize.n431[5] ),
    .B(net699),
    .A(net412));
 sg13g2_or2_1 _3003_ (.X(\serialize.n431[6] ),
    .B(\serialize.n410 ),
    .A(net415));
 sg13g2_mux2_1 _3004_ (.A0(net433),
    .A1(\blue_tmds_par[0] ),
    .S(net699),
    .X(\serialize.n429[0] ));
 sg13g2_mux2_1 _3005_ (.A0(net426),
    .A1(\blue_tmds_par[1] ),
    .S(net699),
    .X(\serialize.n429[1] ));
 sg13g2_mux2_1 _3006_ (.A0(net441),
    .A1(\blue_tmds_par[2] ),
    .S(net695),
    .X(\serialize.n429[2] ));
 sg13g2_mux2_1 _3007_ (.A0(net436),
    .A1(\blue_tmds_par[3] ),
    .S(net695),
    .X(\serialize.n429[3] ));
 sg13g2_mux2_1 _3008_ (.A0(net443),
    .A1(\blue_tmds_par[2] ),
    .S(net695),
    .X(\serialize.n429[4] ));
 sg13g2_mux2_1 _3009_ (.A0(net445),
    .A1(\blue_tmds_par[5] ),
    .S(net695),
    .X(\serialize.n429[5] ));
 sg13g2_mux2_1 _3010_ (.A0(net418),
    .A1(\blue_tmds_par[6] ),
    .S(net695),
    .X(\serialize.n429[6] ));
 sg13g2_mux2_1 _3011_ (.A0(net442),
    .A1(\blue_tmds_par[7] ),
    .S(net696),
    .X(\serialize.n429[7] ));
 sg13g2_and2_1 _3012_ (.A(\blue_tmds_par[8] ),
    .B(net695),
    .X(\serialize.n429[8] ));
 sg13g2_and2_1 _3013_ (.A(\blue_tmds_par[9] ),
    .B(net696),
    .X(\serialize.n429[9] ));
 sg13g2_mux2_1 _3014_ (.A0(net425),
    .A1(\green_tmds_par[0] ),
    .S(net698),
    .X(\serialize.n428[0] ));
 sg13g2_nand2_1 _3015_ (.Y(_0834_),
    .A(\green_tmds_par[1] ),
    .B(net698));
 sg13g2_o21ai_1 _3016_ (.B1(_0834_),
    .Y(\serialize.n428[1] ),
    .A1(_0655_),
    .A2(net700));
 sg13g2_mux2_1 _3017_ (.A0(net440),
    .A1(\green_tmds_par[2] ),
    .S(net697),
    .X(\serialize.n428[2] ));
 sg13g2_o21ai_1 _3018_ (.B1(_0834_),
    .Y(\serialize.n428[3] ),
    .A1(_0656_),
    .A2(net697));
 sg13g2_mux2_1 _3019_ (.A0(net422),
    .A1(\green_tmds_par[2] ),
    .S(net697),
    .X(\serialize.n428[4] ));
 sg13g2_o21ai_1 _3020_ (.B1(_0834_),
    .Y(\serialize.n428[5] ),
    .A1(_0657_),
    .A2(net700));
 sg13g2_mux2_1 _3021_ (.A0(net427),
    .A1(\green_tmds_par[6] ),
    .S(net696),
    .X(\serialize.n428[6] ));
 sg13g2_mux2_1 _3022_ (.A0(net439),
    .A1(\green_tmds_par[7] ),
    .S(net699),
    .X(\serialize.n428[7] ));
 sg13g2_and2_1 _3023_ (.A(\green_tmds_par[8] ),
    .B(net696),
    .X(\serialize.n428[8] ));
 sg13g2_and2_1 _3024_ (.A(\green_tmds_par[9] ),
    .B(net699),
    .X(\serialize.n428[9] ));
 sg13g2_mux2_1 _3025_ (.A0(net438),
    .A1(\red_tmds_par[0] ),
    .S(net698),
    .X(\serialize.n427[0] ));
 sg13g2_mux2_1 _3026_ (.A0(net432),
    .A1(\red_tmds_par[1] ),
    .S(net698),
    .X(\serialize.n427[1] ));
 sg13g2_mux2_1 _3027_ (.A0(net431),
    .A1(\red_tmds_par[2] ),
    .S(net697),
    .X(\serialize.n427[2] ));
 sg13g2_mux2_1 _3028_ (.A0(net437),
    .A1(\red_tmds_par[3] ),
    .S(net697),
    .X(\serialize.n427[3] ));
 sg13g2_mux2_1 _3029_ (.A0(net435),
    .A1(\red_tmds_par[4] ),
    .S(net697),
    .X(\serialize.n427[4] ));
 sg13g2_mux2_1 _3030_ (.A0(net423),
    .A1(\red_tmds_par[5] ),
    .S(net697),
    .X(\serialize.n427[5] ));
 sg13g2_mux2_1 _3031_ (.A0(net419),
    .A1(\red_tmds_par[6] ),
    .S(net696),
    .X(\serialize.n427[6] ));
 sg13g2_mux2_1 _3032_ (.A0(net424),
    .A1(\red_tmds_par[7] ),
    .S(net697),
    .X(\serialize.n427[7] ));
 sg13g2_and2_1 _3033_ (.A(\red_tmds_par[8] ),
    .B(net696),
    .X(\serialize.n427[8] ));
 sg13g2_and2_1 _3034_ (.A(\red_tmds_par[9] ),
    .B(net696),
    .X(\serialize.n427[9] ));
 sg13g2_nor2_1 _3035_ (.A(net679),
    .B(net730),
    .Y(_0006_));
 sg13g2_inv_1 _3036_ (.Y(clk_video),
    .A(_0006_));
 sg13g2_nand2_1 _3037_ (.Y(_0835_),
    .A(net794),
    .B(_0807_));
 sg13g2_nor2_1 _3038_ (.A(_0808_),
    .B(_0835_),
    .Y(_0001_));
 sg13g2_nor2_1 _3039_ (.A(_0807_),
    .B(_0810_),
    .Y(_0000_));
 sg13g2_nor2_2 _3040_ (.A(_0647_),
    .B(net750),
    .Y(_0836_));
 sg13g2_nand2_1 _3041_ (.Y(_0837_),
    .A(net606),
    .B(net796));
 sg13g2_and2_1 _3042_ (.A(\tmds_green.dc_balancing_reg[0] ),
    .B(_0836_),
    .X(_0263_));
 sg13g2_and2_1 _3043_ (.A(\tmds_blue.dc_balancing_reg[0] ),
    .B(_0836_),
    .X(_0264_));
 sg13g2_o21ai_1 _3044_ (.B1(net794),
    .Y(_0838_),
    .A1(net741),
    .A2(net434));
 sg13g2_a21oi_1 _3045_ (.A1(net742),
    .A2(net434),
    .Y(_0265_),
    .B1(_0838_));
 sg13g2_and3_1 _3046_ (.X(_0266_),
    .A(net794),
    .B(net742),
    .C(net434));
 sg13g2_nor2_1 _3047_ (.A(_0642_),
    .B(net569),
    .Y(_0271_));
 sg13g2_nor4_1 _3048_ (.A(\tmds_green.dc_balancing_reg[0] ),
    .B(\tmds_green.dc_balancing_reg[1] ),
    .C(\tmds_green.dc_balancing_reg[3] ),
    .D(\tmds_green.dc_balancing_reg[2] ),
    .Y(_0839_));
 sg13g2_and2_1 _3049_ (.A(_0642_),
    .B(_0839_),
    .X(_0840_));
 sg13g2_nand2b_1 _3050_ (.Y(_0841_),
    .B(net602),
    .A_N(net601));
 sg13g2_xor2_1 _3051_ (.B(net601),
    .A(net602),
    .X(_0842_));
 sg13g2_nand2_1 _3052_ (.Y(_0843_),
    .A(\tmds_green.n100 ),
    .B(_0642_));
 sg13g2_nand2_2 _3053_ (.Y(_0844_),
    .A(net602),
    .B(_0840_));
 sg13g2_mux2_1 _3054_ (.A0(_0842_),
    .A1(net601),
    .S(_0840_),
    .X(_0845_));
 sg13g2_nand2b_1 _3055_ (.Y(_0846_),
    .B(\tmds_green.dc_balancing_reg[4] ),
    .A_N(net603));
 sg13g2_o21ai_1 _3056_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_0839_),
    .A2(_0843_));
 sg13g2_xor2_1 _3057_ (.B(_0847_),
    .A(\tmds_green.n126 ),
    .X(_0848_));
 sg13g2_xnor2_1 _3058_ (.Y(_0849_),
    .A(_0845_),
    .B(_0848_));
 sg13g2_nor2_1 _3059_ (.A(net569),
    .B(_0849_),
    .Y(_0273_));
 sg13g2_a21oi_1 _3060_ (.A1(\tmds_red.n126 ),
    .A2(\tmds_red.n132 ),
    .Y(_0850_),
    .B1(\tmds_red.n102 ));
 sg13g2_nor2_1 _3061_ (.A(\tmds_red.n126 ),
    .B(\tmds_red.n132 ),
    .Y(_0851_));
 sg13g2_nor2_1 _3062_ (.A(\tmds_red.n100 ),
    .B(\tmds_red.n114 ),
    .Y(_0852_));
 sg13g2_nor3_1 _3063_ (.A(_0850_),
    .B(_0851_),
    .C(_0852_),
    .Y(_0853_));
 sg13g2_xnor2_1 _3064_ (.Y(_0854_),
    .A(\tmds_red.n126 ),
    .B(\tmds_red.n132 ));
 sg13g2_a21oi_2 _3065_ (.B1(_0853_),
    .Y(_0855_),
    .A2(\tmds_red.n114 ),
    .A1(\tmds_red.n100 ));
 sg13g2_nor4_1 _3066_ (.A(\tmds_red.dc_balancing_reg[1] ),
    .B(\tmds_red.dc_balancing_reg[0] ),
    .C(\tmds_red.dc_balancing_reg[3] ),
    .D(\tmds_red.dc_balancing_reg[2] ),
    .Y(_0856_));
 sg13g2_nand2_1 _3067_ (.Y(_0857_),
    .A(\tmds_red.n114 ),
    .B(\tmds_red.n132 ));
 sg13g2_nor2_1 _3068_ (.A(\tmds_red.n114 ),
    .B(\tmds_red.n132 ),
    .Y(_0858_));
 sg13g2_xor2_1 _3069_ (.B(\tmds_red.n132 ),
    .A(\tmds_red.n114 ),
    .X(_0859_));
 sg13g2_xnor2_1 _3070_ (.Y(_0860_),
    .A(\tmds_red.n100 ),
    .B(\tmds_red.n102 ));
 sg13g2_xnor2_1 _3071_ (.Y(_0861_),
    .A(net548),
    .B(_0860_));
 sg13g2_xnor2_1 _3072_ (.Y(_0862_),
    .A(_0859_),
    .B(_0861_));
 sg13g2_nor2_1 _3073_ (.A(\tmds_red.n102 ),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_nand2_1 _3074_ (.Y(_0864_),
    .A(\tmds_red.n102 ),
    .B(_0862_));
 sg13g2_nand2b_1 _3075_ (.Y(_0865_),
    .B(\tmds_red.n100 ),
    .A_N(_0859_));
 sg13g2_a21oi_1 _3076_ (.A1(_0857_),
    .A2(_0860_),
    .Y(_0866_),
    .B1(_0858_));
 sg13g2_nor2b_1 _3077_ (.A(\tmds_red.n126 ),
    .B_N(\tmds_red.n132 ),
    .Y(_0867_));
 sg13g2_a21oi_1 _3078_ (.A1(_0854_),
    .A2(net548),
    .Y(_0868_),
    .B1(_0867_));
 sg13g2_xnor2_1 _3079_ (.Y(_0869_),
    .A(_0866_),
    .B(_0868_));
 sg13g2_nand2_1 _3080_ (.Y(_0870_),
    .A(_0861_),
    .B(_0869_));
 sg13g2_xnor2_1 _3081_ (.Y(_0871_),
    .A(_0859_),
    .B(_0869_));
 sg13g2_nor2_1 _3082_ (.A(_0861_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_a21o_1 _3083_ (.A2(_0869_),
    .A1(_0861_),
    .B1(_0872_),
    .X(_0873_));
 sg13g2_o21ai_1 _3084_ (.B1(_0864_),
    .Y(_0874_),
    .A1(net548),
    .A2(_0863_));
 sg13g2_xnor2_1 _3085_ (.Y(_0875_),
    .A(_0873_),
    .B(_0874_));
 sg13g2_nor2b_1 _3086_ (.A(_0865_),
    .B_N(_0875_),
    .Y(_0876_));
 sg13g2_o21ai_1 _3087_ (.B1(_0870_),
    .Y(_0877_),
    .A1(_0872_),
    .A2(_0874_));
 sg13g2_nor2b_2 _3088_ (.A(_0877_),
    .B_N(_0876_),
    .Y(_0878_));
 sg13g2_nand2b_1 _3089_ (.Y(_0879_),
    .B(_0877_),
    .A_N(_0876_));
 sg13g2_inv_2 _3090_ (.Y(_0880_),
    .A(_0879_));
 sg13g2_nor2_1 _3091_ (.A(_0878_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_xnor2_1 _3092_ (.Y(_0882_),
    .A(_0865_),
    .B(_0875_));
 sg13g2_nor2_2 _3093_ (.A(_0859_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_a22oi_1 _3094_ (.Y(_0884_),
    .B1(_0881_),
    .B2(_0883_),
    .A2(_0856_),
    .A1(_0652_));
 sg13g2_nor2b_2 _3095_ (.A(_0884_),
    .B_N(net548),
    .Y(_0885_));
 sg13g2_nor3_1 _3096_ (.A(_0878_),
    .B(_0880_),
    .C(_0883_),
    .Y(_0886_));
 sg13g2_nor2_1 _3097_ (.A(_0878_),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_nor3_1 _3098_ (.A(\tmds_red.dc_balancing_reg[4] ),
    .B(_0856_),
    .C(_0887_),
    .Y(_0888_));
 sg13g2_a21oi_2 _3099_ (.B1(_0888_),
    .Y(_0889_),
    .A2(_0880_),
    .A1(\tmds_red.dc_balancing_reg[4] ));
 sg13g2_nand2_1 _3100_ (.Y(_0890_),
    .A(_0884_),
    .B(_0889_));
 sg13g2_a21oi_2 _3101_ (.B1(_0885_),
    .Y(_0891_),
    .A2(_0889_),
    .A1(_0884_));
 sg13g2_o21ai_1 _3102_ (.B1(_0836_),
    .Y(_0892_),
    .A1(\tmds_red.n100 ),
    .A2(_0891_));
 sg13g2_a21oi_1 _3103_ (.A1(\tmds_red.n100 ),
    .A2(_0891_),
    .Y(_0274_),
    .B1(_0892_));
 sg13g2_mux2_1 _3104_ (.A0(_0890_),
    .A1(_0889_),
    .S(net548),
    .X(_0893_));
 sg13g2_nor2_1 _3105_ (.A(net570),
    .B(_0893_),
    .Y(_0275_));
 sg13g2_xnor2_1 _3106_ (.Y(_0894_),
    .A(_0860_),
    .B(_0893_));
 sg13g2_nor2_1 _3107_ (.A(net569),
    .B(_0894_),
    .Y(_0276_));
 sg13g2_xnor2_1 _3108_ (.Y(_0895_),
    .A(_0854_),
    .B(_0894_));
 sg13g2_nor2_1 _3109_ (.A(net569),
    .B(_0895_),
    .Y(_0278_));
 sg13g2_nor3_1 _3110_ (.A(net629),
    .B(\videogen.fancy_shader.video_x[6] ),
    .C(\videogen.fancy_shader.video_x[5] ),
    .Y(_0896_));
 sg13g2_and3_2 _3111_ (.X(_0897_),
    .A(_0791_),
    .B(_0798_),
    .C(_0896_));
 sg13g2_nand2b_2 _3112_ (.Y(_0898_),
    .B(net795),
    .A_N(_0897_));
 sg13g2_nor2_1 _3113_ (.A(net630),
    .B(_0898_),
    .Y(_0303_));
 sg13g2_xnor2_1 _3114_ (.Y(_0899_),
    .A(\videogen.fancy_shader.video_x[1] ),
    .B(net630));
 sg13g2_nor2_1 _3115_ (.A(_0898_),
    .B(_0899_),
    .Y(_0304_));
 sg13g2_a21oi_1 _3116_ (.A1(\videogen.fancy_shader.video_x[1] ),
    .A2(net630),
    .Y(_0900_),
    .B1(\videogen.fancy_shader.video_x[2] ));
 sg13g2_nor3_1 _3117_ (.A(net751),
    .B(_0795_),
    .C(_0900_),
    .Y(_0305_));
 sg13g2_o21ai_1 _3118_ (.B1(net795),
    .Y(_0901_),
    .A1(\videogen.fancy_shader.video_x[3] ),
    .A2(_0795_));
 sg13g2_nor2_1 _3119_ (.A(_0796_),
    .B(_0901_),
    .Y(_0306_));
 sg13g2_nand2b_1 _3120_ (.Y(_0902_),
    .B(_0797_),
    .A_N(\videogen.fancy_shader.video_x[4] ));
 sg13g2_nand2_1 _3121_ (.Y(_0903_),
    .A(net795),
    .B(_0902_));
 sg13g2_nor2_1 _3122_ (.A(_0798_),
    .B(_0903_),
    .Y(_0307_));
 sg13g2_nor2_1 _3123_ (.A(\videogen.fancy_shader.video_x[5] ),
    .B(_0798_),
    .Y(_0904_));
 sg13g2_nor3_1 _3124_ (.A(_0799_),
    .B(_0898_),
    .C(_0904_),
    .Y(_0308_));
 sg13g2_nor2_1 _3125_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(_0799_),
    .Y(_0905_));
 sg13g2_nor3_1 _3126_ (.A(_0800_),
    .B(_0898_),
    .C(_0905_),
    .Y(_0309_));
 sg13g2_and2_1 _3127_ (.A(net629),
    .B(_0800_),
    .X(_0906_));
 sg13g2_nor2_1 _3128_ (.A(net629),
    .B(_0800_),
    .Y(_0907_));
 sg13g2_nor3_1 _3129_ (.A(_0898_),
    .B(_0906_),
    .C(_0907_),
    .Y(_0310_));
 sg13g2_nand2_1 _3130_ (.Y(_0908_),
    .A(\videogen.fancy_shader.video_x[8] ),
    .B(_0906_));
 sg13g2_xnor2_1 _3131_ (.Y(_0909_),
    .A(\videogen.fancy_shader.video_x[8] ),
    .B(_0906_));
 sg13g2_nor2_1 _3132_ (.A(_0898_),
    .B(_0909_),
    .Y(_0311_));
 sg13g2_xor2_1 _3133_ (.B(_0908_),
    .A(\videogen.fancy_shader.video_x[9] ),
    .X(_0910_));
 sg13g2_nor2_1 _3134_ (.A(_0898_),
    .B(_0910_),
    .Y(_0312_));
 sg13g2_nand2b_1 _3135_ (.Y(_0911_),
    .B(\videogen.fancy_shader.video_y[3] ),
    .A_N(\videogen.fancy_shader.video_y[2] ));
 sg13g2_nor4_1 _3136_ (.A(_0662_),
    .B(_0663_),
    .C(_0814_),
    .D(_0911_),
    .Y(_0912_));
 sg13g2_nor2_1 _3137_ (.A(net748),
    .B(_0912_),
    .Y(_0317_));
 sg13g2_nor3_1 _3138_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .Y(_0913_));
 sg13g2_o21ai_1 _3139_ (.B1(_0672_),
    .Y(_0914_),
    .A1(\videogen.mem_read ),
    .A2(_0809_));
 sg13g2_nor2b_1 _3140_ (.A(_0914_),
    .B_N(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .Y(_0915_));
 sg13g2_nor2b_1 _3141_ (.A(_0913_),
    .B_N(_0915_),
    .Y(_0916_));
 sg13g2_nor2_1 _3142_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nand2_2 _3143_ (.Y(_0918_),
    .A(_0665_),
    .B(_0670_));
 sg13g2_nand2_2 _3144_ (.Y(_0919_),
    .A(net793),
    .B(_0918_));
 sg13g2_and2_1 _3145_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0916_),
    .X(_0920_));
 sg13g2_nor3_1 _3146_ (.A(_0917_),
    .B(_0919_),
    .C(_0920_),
    .Y(_0318_));
 sg13g2_nor2_1 _3147_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_and2_1 _3148_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .B(_0920_),
    .X(_0922_));
 sg13g2_nor3_1 _3149_ (.A(_0919_),
    .B(_0921_),
    .C(_0922_),
    .Y(_0319_));
 sg13g2_and2_1 _3150_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(_0922_),
    .X(_0923_));
 sg13g2_nor2_1 _3151_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(_0922_),
    .Y(_0924_));
 sg13g2_nor3_1 _3152_ (.A(_0919_),
    .B(_0923_),
    .C(_0924_),
    .Y(_0320_));
 sg13g2_and2_1 _3153_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B(_0923_),
    .X(_0925_));
 sg13g2_nor2_1 _3154_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B(_0923_),
    .Y(_0926_));
 sg13g2_nor3_1 _3155_ (.A(_0919_),
    .B(_0925_),
    .C(_0926_),
    .Y(_0321_));
 sg13g2_nor2_1 _3156_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .B(_0925_),
    .Y(_0927_));
 sg13g2_and2_1 _3157_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .B(_0925_),
    .X(_0928_));
 sg13g2_nor3_1 _3158_ (.A(_0919_),
    .B(_0927_),
    .C(_0928_),
    .Y(_0322_));
 sg13g2_a21oi_1 _3159_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0928_),
    .Y(_0929_),
    .B1(_0919_));
 sg13g2_o21ai_1 _3160_ (.B1(_0929_),
    .Y(_0930_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0928_));
 sg13g2_inv_1 _3161_ (.Y(_0323_),
    .A(_0930_));
 sg13g2_nor3_1 _3162_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .Y(_0931_));
 sg13g2_nand2_1 _3163_ (.Y(_0932_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .B(_0792_));
 sg13g2_nor2_1 _3164_ (.A(_0931_),
    .B(_0932_),
    .Y(_0933_));
 sg13g2_xnor2_1 _3165_ (.Y(_0934_),
    .A(net628),
    .B(_0933_));
 sg13g2_nor2_1 _3166_ (.A(_0793_),
    .B(_0934_),
    .Y(_0324_));
 sg13g2_nor3_1 _3167_ (.A(net578),
    .B(_0931_),
    .C(_0932_),
    .Y(_0935_));
 sg13g2_a21oi_1 _3168_ (.A1(net628),
    .A2(_0933_),
    .Y(_0936_),
    .B1(net625));
 sg13g2_nor3_1 _3169_ (.A(_0793_),
    .B(_0935_),
    .C(_0936_),
    .Y(_0325_));
 sg13g2_nor2_1 _3170_ (.A(net621),
    .B(_0935_),
    .Y(_0937_));
 sg13g2_and2_1 _3171_ (.A(net621),
    .B(_0935_),
    .X(_0938_));
 sg13g2_nor3_1 _3172_ (.A(_0793_),
    .B(_0937_),
    .C(_0938_),
    .Y(_0326_));
 sg13g2_xnor2_1 _3173_ (.Y(_0939_),
    .A(net616),
    .B(_0938_));
 sg13g2_nor2_1 _3174_ (.A(_0793_),
    .B(_0939_),
    .Y(_0327_));
 sg13g2_a21oi_1 _3175_ (.A1(net616),
    .A2(_0938_),
    .Y(_0940_),
    .B1(net613));
 sg13g2_nand3_1 _3176_ (.B(net616),
    .C(_0938_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .Y(_0941_));
 sg13g2_nand2_1 _3177_ (.Y(_0942_),
    .A(_0794_),
    .B(_0941_));
 sg13g2_nor2_1 _3178_ (.A(_0940_),
    .B(_0942_),
    .Y(_0328_));
 sg13g2_xnor2_1 _3179_ (.Y(_0943_),
    .A(_0636_),
    .B(_0941_));
 sg13g2_nor2_1 _3180_ (.A(_0793_),
    .B(_0943_),
    .Y(_0329_));
 sg13g2_or2_1 _3181_ (.X(_0944_),
    .B(_0919_),
    .A(_0916_));
 sg13g2_nor2b_1 _3182_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .B_N(_0914_),
    .Y(_0945_));
 sg13g2_nor2b_1 _3183_ (.A(_0914_),
    .B_N(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .Y(_0946_));
 sg13g2_nor3_1 _3184_ (.A(_0944_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0330_));
 sg13g2_nor2_1 _3185_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_and2_1 _3186_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .B(_0946_),
    .X(_0948_));
 sg13g2_nor4_1 _3187_ (.A(_0915_),
    .B(_0919_),
    .C(_0947_),
    .D(_0948_),
    .Y(_0331_));
 sg13g2_xnor2_1 _3188_ (.Y(_0949_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .B(_0948_));
 sg13g2_nor2_1 _3189_ (.A(_0944_),
    .B(_0949_),
    .Y(_0332_));
 sg13g2_a21oi_1 _3190_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .A2(_0948_),
    .Y(_0950_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ));
 sg13g2_nor2_1 _3191_ (.A(_0944_),
    .B(_0950_),
    .Y(_0333_));
 sg13g2_o21ai_1 _3192_ (.B1(_0794_),
    .Y(_0951_),
    .A1(_0931_),
    .A2(_0932_));
 sg13g2_nor2_1 _3193_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .B(_0792_),
    .Y(_0952_));
 sg13g2_nor3_1 _3194_ (.A(_0802_),
    .B(_0951_),
    .C(_0952_),
    .Y(_0334_));
 sg13g2_nor2_1 _3195_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .B(_0802_),
    .Y(_0953_));
 sg13g2_and2_1 _3196_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .B(_0802_),
    .X(_0954_));
 sg13g2_nor3_1 _3197_ (.A(_0951_),
    .B(_0953_),
    .C(_0954_),
    .Y(_0335_));
 sg13g2_xnor2_1 _3198_ (.Y(_0955_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(_0954_));
 sg13g2_nor2_1 _3199_ (.A(_0951_),
    .B(_0955_),
    .Y(_0336_));
 sg13g2_a21oi_1 _3200_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .A2(_0954_),
    .Y(_0956_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ));
 sg13g2_nor2_1 _3201_ (.A(_0951_),
    .B(_0956_),
    .Y(_0337_));
 sg13g2_nor2_1 _3202_ (.A(_0635_),
    .B(_0918_),
    .Y(_0957_));
 sg13g2_a21oi_1 _3203_ (.A1(_0635_),
    .A2(_0918_),
    .Y(_0958_),
    .B1(net751));
 sg13g2_nor2b_1 _3204_ (.A(_0957_),
    .B_N(_0958_),
    .Y(_0346_));
 sg13g2_nor2_1 _3205_ (.A(\videogen.fancy_shader.n646[1] ),
    .B(_0957_),
    .Y(_0959_));
 sg13g2_and2_1 _3206_ (.A(\videogen.fancy_shader.n646[1] ),
    .B(_0957_),
    .X(_0960_));
 sg13g2_nor3_1 _3207_ (.A(net751),
    .B(_0959_),
    .C(_0960_),
    .Y(_0347_));
 sg13g2_and2_1 _3208_ (.A(\videogen.fancy_shader.n646[2] ),
    .B(_0960_),
    .X(_0961_));
 sg13g2_o21ai_1 _3209_ (.B1(net795),
    .Y(_0962_),
    .A1(\videogen.fancy_shader.n646[2] ),
    .A2(_0960_));
 sg13g2_nor2_1 _3210_ (.A(_0961_),
    .B(_0962_),
    .Y(_0348_));
 sg13g2_xnor2_1 _3211_ (.Y(_0963_),
    .A(\videogen.fancy_shader.n646[3] ),
    .B(_0961_));
 sg13g2_nor2_1 _3212_ (.A(net751),
    .B(_0963_),
    .Y(_0349_));
 sg13g2_a21oi_1 _3213_ (.A1(net611),
    .A2(_0961_),
    .Y(_0964_),
    .B1(\videogen.fancy_shader.n646[4] ));
 sg13g2_and3_2 _3214_ (.X(_0965_),
    .A(\videogen.fancy_shader.n646[4] ),
    .B(net611),
    .C(_0961_));
 sg13g2_nor3_1 _3215_ (.A(net751),
    .B(_0964_),
    .C(_0965_),
    .Y(_0350_));
 sg13g2_xnor2_1 _3216_ (.Y(_0966_),
    .A(\videogen.fancy_shader.n646[5] ),
    .B(_0965_));
 sg13g2_nor2_1 _3217_ (.A(net747),
    .B(_0966_),
    .Y(_0351_));
 sg13g2_a21oi_1 _3218_ (.A1(\videogen.fancy_shader.n646[5] ),
    .A2(_0965_),
    .Y(_0967_),
    .B1(\videogen.fancy_shader.n646[6] ));
 sg13g2_and3_1 _3219_ (.X(_0968_),
    .A(\videogen.fancy_shader.n646[6] ),
    .B(\videogen.fancy_shader.n646[5] ),
    .C(_0965_));
 sg13g2_nor3_1 _3220_ (.A(net748),
    .B(_0967_),
    .C(_0968_),
    .Y(_0352_));
 sg13g2_nor2_1 _3221_ (.A(\videogen.fancy_shader.n646[7] ),
    .B(_0968_),
    .Y(_0969_));
 sg13g2_and2_1 _3222_ (.A(\videogen.fancy_shader.n646[7] ),
    .B(_0968_),
    .X(_0970_));
 sg13g2_nor3_1 _3223_ (.A(net747),
    .B(_0969_),
    .C(_0970_),
    .Y(_0353_));
 sg13g2_xnor2_1 _3224_ (.Y(_0971_),
    .A(net610),
    .B(_0970_));
 sg13g2_nor2_1 _3225_ (.A(net747),
    .B(_0971_),
    .Y(_0354_));
 sg13g2_a21oi_1 _3226_ (.A1(net610),
    .A2(_0970_),
    .Y(_0972_),
    .B1(\videogen.fancy_shader.n646[9] ));
 sg13g2_and3_1 _3227_ (.X(_0973_),
    .A(\videogen.fancy_shader.n646[9] ),
    .B(\videogen.fancy_shader.n646[8] ),
    .C(_0970_));
 sg13g2_nor3_1 _3228_ (.A(net747),
    .B(_0972_),
    .C(_0973_),
    .Y(_0355_));
 sg13g2_and2_1 _3229_ (.A(net609),
    .B(_0897_),
    .X(_0974_));
 sg13g2_o21ai_1 _3230_ (.B1(net795),
    .Y(_0975_),
    .A1(net609),
    .A2(_0897_));
 sg13g2_nor2_1 _3231_ (.A(_0974_),
    .B(_0975_),
    .Y(_0356_));
 sg13g2_and2_1 _3232_ (.A(net608),
    .B(_0974_),
    .X(_0976_));
 sg13g2_o21ai_1 _3233_ (.B1(net803),
    .Y(_0977_),
    .A1(net608),
    .A2(_0974_));
 sg13g2_nor2_1 _3234_ (.A(_0976_),
    .B(_0977_),
    .Y(_0357_));
 sg13g2_nor4_1 _3235_ (.A(\videogen.fancy_shader.video_y[7] ),
    .B(\videogen.fancy_shader.video_y[6] ),
    .C(\videogen.fancy_shader.video_y[5] ),
    .D(\videogen.fancy_shader.video_y[4] ),
    .Y(_0978_));
 sg13g2_nor4_1 _3236_ (.A(_0632_),
    .B(\videogen.fancy_shader.video_y[8] ),
    .C(_0815_),
    .D(_0911_),
    .Y(_0979_));
 sg13g2_nand3_1 _3237_ (.B(_0978_),
    .C(_0979_),
    .A(_0897_),
    .Y(_0980_));
 sg13g2_nand2_1 _3238_ (.Y(_0981_),
    .A(net795),
    .B(_0980_));
 sg13g2_xnor2_1 _3239_ (.Y(_0982_),
    .A(\videogen.fancy_shader.video_y[2] ),
    .B(_0976_));
 sg13g2_nor2_1 _3240_ (.A(_0981_),
    .B(_0982_),
    .Y(_0358_));
 sg13g2_a22oi_1 _3241_ (.Y(_0983_),
    .B1(_0980_),
    .B2(\videogen.fancy_shader.video_y[3] ),
    .A2(_0976_),
    .A1(\videogen.fancy_shader.video_y[2] ));
 sg13g2_and4_1 _3242_ (.A(\videogen.fancy_shader.video_y[3] ),
    .B(\videogen.fancy_shader.video_y[2] ),
    .C(_0814_),
    .D(_0897_),
    .X(_0984_));
 sg13g2_nor3_1 _3243_ (.A(net748),
    .B(_0983_),
    .C(_0984_),
    .Y(_0359_));
 sg13g2_nor2b_1 _3244_ (.A(_0816_),
    .B_N(_0976_),
    .Y(_0985_));
 sg13g2_o21ai_1 _3245_ (.B1(net795),
    .Y(_0986_),
    .A1(\videogen.fancy_shader.video_y[4] ),
    .A2(_0984_));
 sg13g2_nor2_1 _3246_ (.A(_0985_),
    .B(_0986_),
    .Y(_0360_));
 sg13g2_nor2_1 _3247_ (.A(\videogen.fancy_shader.video_y[5] ),
    .B(_0985_),
    .Y(_0987_));
 sg13g2_and3_2 _3248_ (.X(_0988_),
    .A(\videogen.fancy_shader.video_y[5] ),
    .B(\videogen.fancy_shader.video_y[4] ),
    .C(_0984_));
 sg13g2_nor3_1 _3249_ (.A(net748),
    .B(_0987_),
    .C(_0988_),
    .Y(_0361_));
 sg13g2_xnor2_1 _3250_ (.Y(_0989_),
    .A(\videogen.fancy_shader.video_y[6] ),
    .B(_0988_));
 sg13g2_nor2_1 _3251_ (.A(net747),
    .B(_0989_),
    .Y(_0362_));
 sg13g2_a21oi_1 _3252_ (.A1(\videogen.fancy_shader.video_y[6] ),
    .A2(_0988_),
    .Y(_0990_),
    .B1(\videogen.fancy_shader.video_y[7] ));
 sg13g2_and3_1 _3253_ (.X(_0991_),
    .A(\videogen.fancy_shader.video_y[7] ),
    .B(\videogen.fancy_shader.video_y[6] ),
    .C(_0988_));
 sg13g2_nor3_1 _3254_ (.A(net747),
    .B(_0990_),
    .C(_0991_),
    .Y(_0363_));
 sg13g2_nor2_1 _3255_ (.A(\videogen.fancy_shader.video_y[8] ),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_and2_1 _3256_ (.A(\videogen.fancy_shader.video_y[8] ),
    .B(_0991_),
    .X(_0993_));
 sg13g2_nor3_1 _3257_ (.A(net747),
    .B(_0992_),
    .C(_0993_),
    .Y(_0364_));
 sg13g2_nor2_1 _3258_ (.A(\videogen.fancy_shader.video_y[9] ),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_a21oi_1 _3259_ (.A1(\videogen.fancy_shader.video_y[9] ),
    .A2(_0993_),
    .Y(_0995_),
    .B1(_0981_));
 sg13g2_nor2b_1 _3260_ (.A(_0994_),
    .B_N(_0995_),
    .Y(_0365_));
 sg13g2_nor2_1 _3261_ (.A(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .B(net749),
    .Y(_0366_));
 sg13g2_o21ai_1 _3262_ (.B1(net793),
    .Y(_0996_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ));
 sg13g2_a21oi_1 _3263_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .Y(_0367_),
    .B1(_0996_));
 sg13g2_a21oi_1 _3264_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .Y(_0997_),
    .B1(\videogen.test_lut_thingy.gol_counter_reg[2] ));
 sg13g2_and3_1 _3265_ (.X(_0998_),
    .A(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .B(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .C(\videogen.test_lut_thingy.gol_counter_reg[2] ));
 sg13g2_nor3_1 _3266_ (.A(net749),
    .B(_0997_),
    .C(_0998_),
    .Y(_0368_));
 sg13g2_o21ai_1 _3267_ (.B1(net793),
    .Y(_0999_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A2(_0998_));
 sg13g2_a21oi_1 _3268_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A2(_0998_),
    .Y(_0369_),
    .B1(_0999_));
 sg13g2_nand4_1 _3269_ (.B(\videogen.fancy_shader.video_x[6] ),
    .C(\videogen.fancy_shader.video_x[5] ),
    .A(\videogen.fancy_shader.video_x[7] ),
    .Y(_1000_),
    .D(_0902_));
 sg13g2_nand2_1 _3270_ (.Y(_1001_),
    .A(_0667_),
    .B(_1000_));
 sg13g2_a21oi_1 _3271_ (.A1(_0668_),
    .A2(_0797_),
    .Y(_1002_),
    .B1(_1001_));
 sg13g2_nor2_1 _3272_ (.A(net748),
    .B(_1002_),
    .Y(_0370_));
 sg13g2_nand2_1 _3273_ (.Y(_1003_),
    .A(net608),
    .B(\videogen.fancy_shader.n646[1] ));
 sg13g2_nand2_1 _3274_ (.Y(_1004_),
    .A(net609),
    .B(\videogen.fancy_shader.n646[0] ));
 sg13g2_nor2_1 _3275_ (.A(net608),
    .B(\videogen.fancy_shader.n646[1] ),
    .Y(_1005_));
 sg13g2_xor2_1 _3276_ (.B(\videogen.fancy_shader.n646[1] ),
    .A(\videogen.fancy_shader.video_y[1] ),
    .X(_1006_));
 sg13g2_o21ai_1 _3277_ (.B1(_1003_),
    .Y(_1007_),
    .A1(_1004_),
    .A2(_1005_));
 sg13g2_and2_1 _3278_ (.A(\videogen.fancy_shader.video_y[2] ),
    .B(\videogen.fancy_shader.n646[2] ),
    .X(_1008_));
 sg13g2_xor2_1 _3279_ (.B(\videogen.fancy_shader.n646[2] ),
    .A(\videogen.fancy_shader.video_y[2] ),
    .X(_1009_));
 sg13g2_xnor2_1 _3280_ (.Y(_1010_),
    .A(_1007_),
    .B(_1009_));
 sg13g2_nand2_1 _3281_ (.Y(_1011_),
    .A(\videogen.fancy_shader.n646[1] ),
    .B(\videogen.fancy_shader.video_x[1] ));
 sg13g2_nand2_1 _3282_ (.Y(_1012_),
    .A(\videogen.fancy_shader.n646[0] ),
    .B(net630));
 sg13g2_xnor2_1 _3283_ (.Y(_1013_),
    .A(\videogen.fancy_shader.n646[1] ),
    .B(\videogen.fancy_shader.video_x[1] ));
 sg13g2_o21ai_1 _3284_ (.B1(_1011_),
    .Y(_1014_),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_nand2_1 _3285_ (.Y(_1015_),
    .A(\videogen.fancy_shader.n646[2] ),
    .B(\videogen.fancy_shader.video_x[2] ));
 sg13g2_xnor2_1 _3286_ (.Y(_1016_),
    .A(\videogen.fancy_shader.n646[2] ),
    .B(\videogen.fancy_shader.video_x[2] ));
 sg13g2_nand2b_1 _3287_ (.Y(_1017_),
    .B(_1014_),
    .A_N(_1016_));
 sg13g2_xor2_1 _3288_ (.B(_1016_),
    .A(_1014_),
    .X(_1018_));
 sg13g2_nand2_1 _3289_ (.Y(_1019_),
    .A(_1010_),
    .B(_1018_));
 sg13g2_or2_1 _3290_ (.X(_1020_),
    .B(_1018_),
    .A(_1010_));
 sg13g2_and2_1 _3291_ (.A(_1019_),
    .B(_1020_),
    .X(_1021_));
 sg13g2_inv_1 _3292_ (.Y(_1022_),
    .A(net545));
 sg13g2_nand2_1 _3293_ (.Y(_1023_),
    .A(net611),
    .B(\videogen.fancy_shader.video_x[3] ));
 sg13g2_nor2_1 _3294_ (.A(net611),
    .B(\videogen.fancy_shader.video_x[3] ),
    .Y(_1024_));
 sg13g2_xor2_1 _3295_ (.B(\videogen.fancy_shader.video_x[3] ),
    .A(net611),
    .X(_1025_));
 sg13g2_and2_1 _3296_ (.A(_1015_),
    .B(_1017_),
    .X(_1026_));
 sg13g2_xnor2_1 _3297_ (.Y(_1027_),
    .A(_1025_),
    .B(_1026_));
 sg13g2_nor2_1 _3298_ (.A(\videogen.fancy_shader.video_y[3] ),
    .B(net611),
    .Y(_1028_));
 sg13g2_xor2_1 _3299_ (.B(net611),
    .A(\videogen.fancy_shader.video_y[3] ),
    .X(_1029_));
 sg13g2_a21oi_1 _3300_ (.A1(_1007_),
    .A2(_1009_),
    .Y(_1030_),
    .B1(_1008_));
 sg13g2_xnor2_1 _3301_ (.Y(_1031_),
    .A(_1029_),
    .B(_1030_));
 sg13g2_or2_1 _3302_ (.X(_1032_),
    .B(net546),
    .A(_1027_));
 sg13g2_nand2_1 _3303_ (.Y(_1033_),
    .A(_1027_),
    .B(net546));
 sg13g2_nand2b_1 _3304_ (.Y(_1034_),
    .B(_1027_),
    .A_N(net546));
 sg13g2_nand2b_1 _3305_ (.Y(_1035_),
    .B(net546),
    .A_N(_1027_));
 sg13g2_nand2_2 _3306_ (.Y(_1036_),
    .A(_1034_),
    .B(_1035_));
 sg13g2_inv_1 _3307_ (.Y(_1037_),
    .A(_1036_));
 sg13g2_nor2b_1 _3308_ (.A(_1016_),
    .B_N(_1025_),
    .Y(_1038_));
 sg13g2_inv_1 _3309_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_o21ai_1 _3310_ (.B1(_1023_),
    .Y(_1040_),
    .A1(_1015_),
    .A2(_1024_));
 sg13g2_a21oi_1 _3311_ (.A1(_1014_),
    .A2(_1038_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_a21o_1 _3312_ (.A2(_1038_),
    .A1(_1014_),
    .B1(_1040_),
    .X(_1042_));
 sg13g2_nand2_1 _3313_ (.Y(_1043_),
    .A(\videogen.fancy_shader.n646[4] ),
    .B(\videogen.fancy_shader.video_x[4] ));
 sg13g2_xor2_1 _3314_ (.B(\videogen.fancy_shader.video_x[4] ),
    .A(\videogen.fancy_shader.n646[4] ),
    .X(_1044_));
 sg13g2_nand2_1 _3315_ (.Y(_1045_),
    .A(_1042_),
    .B(_1044_));
 sg13g2_xnor2_1 _3316_ (.Y(_1046_),
    .A(_1041_),
    .B(_1044_));
 sg13g2_and2_1 _3317_ (.A(_1009_),
    .B(_1029_),
    .X(_1047_));
 sg13g2_nor2b_1 _3318_ (.A(_1028_),
    .B_N(_1008_),
    .Y(_1048_));
 sg13g2_a221oi_1 _3319_ (.B2(_1047_),
    .C1(_1048_),
    .B1(_1007_),
    .A1(\videogen.fancy_shader.video_y[3] ),
    .Y(_1049_),
    .A2(net611));
 sg13g2_nand2_1 _3320_ (.Y(_1050_),
    .A(\videogen.fancy_shader.video_y[4] ),
    .B(\videogen.fancy_shader.n646[4] ));
 sg13g2_xnor2_1 _3321_ (.Y(_1051_),
    .A(\videogen.fancy_shader.video_y[4] ),
    .B(\videogen.fancy_shader.n646[4] ));
 sg13g2_xor2_1 _3322_ (.B(_1051_),
    .A(_1049_),
    .X(_1052_));
 sg13g2_or2_1 _3323_ (.X(_1053_),
    .B(_1052_),
    .A(_1046_));
 sg13g2_nand2_1 _3324_ (.Y(_1054_),
    .A(_1046_),
    .B(_1052_));
 sg13g2_nand2_2 _3325_ (.Y(_1055_),
    .A(_1053_),
    .B(_1054_));
 sg13g2_inv_1 _3326_ (.Y(_1056_),
    .A(net544));
 sg13g2_nand2_1 _3327_ (.Y(_1057_),
    .A(_0634_),
    .B(_0640_));
 sg13g2_xor2_1 _3328_ (.B(\videogen.fancy_shader.video_x[5] ),
    .A(\videogen.fancy_shader.n646[5] ),
    .X(_1058_));
 sg13g2_nand2_1 _3329_ (.Y(_1059_),
    .A(_1043_),
    .B(_1045_));
 sg13g2_xnor2_1 _3330_ (.Y(_1060_),
    .A(_1058_),
    .B(_1059_));
 sg13g2_xnor2_1 _3331_ (.Y(_1061_),
    .A(\videogen.fancy_shader.video_y[5] ),
    .B(\videogen.fancy_shader.n646[5] ));
 sg13g2_o21ai_1 _3332_ (.B1(_1050_),
    .Y(_1062_),
    .A1(_1049_),
    .A2(_1051_));
 sg13g2_xnor2_1 _3333_ (.Y(_1063_),
    .A(_1061_),
    .B(_1062_));
 sg13g2_or2_1 _3334_ (.X(_1064_),
    .B(_1063_),
    .A(_1060_));
 sg13g2_nand2_1 _3335_ (.Y(_1065_),
    .A(_1060_),
    .B(_1063_));
 sg13g2_and2_1 _3336_ (.A(_1064_),
    .B(_1065_),
    .X(_1066_));
 sg13g2_inv_1 _3337_ (.Y(_1067_),
    .A(_1066_));
 sg13g2_nand2_1 _3338_ (.Y(_1068_),
    .A(_1044_),
    .B(_1058_));
 sg13g2_inv_1 _3339_ (.Y(_1069_),
    .A(_1068_));
 sg13g2_o21ai_1 _3340_ (.B1(_1043_),
    .Y(_1070_),
    .A1(_0634_),
    .A2(_0640_));
 sg13g2_nand2_1 _3341_ (.Y(_1071_),
    .A(_1057_),
    .B(_1070_));
 sg13g2_a22oi_1 _3342_ (.Y(_1072_),
    .B1(_1070_),
    .B2(_1057_),
    .A2(_1069_),
    .A1(_1042_));
 sg13g2_o21ai_1 _3343_ (.B1(_1071_),
    .Y(_1073_),
    .A1(_1041_),
    .A2(_1068_));
 sg13g2_nand2_1 _3344_ (.Y(_1074_),
    .A(\videogen.fancy_shader.n646[6] ),
    .B(\videogen.fancy_shader.video_x[6] ));
 sg13g2_xnor2_1 _3345_ (.Y(_1075_),
    .A(\videogen.fancy_shader.n646[6] ),
    .B(\videogen.fancy_shader.video_x[6] ));
 sg13g2_xnor2_1 _3346_ (.Y(_1076_),
    .A(_1073_),
    .B(_1075_));
 sg13g2_or2_1 _3347_ (.X(_1077_),
    .B(_1061_),
    .A(_1051_));
 sg13g2_o21ai_1 _3348_ (.B1(_1050_),
    .Y(_1078_),
    .A1(_0633_),
    .A2(_0634_));
 sg13g2_o21ai_1 _3349_ (.B1(_1078_),
    .Y(_1079_),
    .A1(\videogen.fancy_shader.video_y[5] ),
    .A2(\videogen.fancy_shader.n646[5] ));
 sg13g2_o21ai_1 _3350_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1049_),
    .A2(_1077_));
 sg13g2_and2_1 _3351_ (.A(\videogen.fancy_shader.video_y[6] ),
    .B(\videogen.fancy_shader.n646[6] ),
    .X(_1081_));
 sg13g2_or2_1 _3352_ (.X(_1082_),
    .B(\videogen.fancy_shader.n646[6] ),
    .A(\videogen.fancy_shader.video_y[6] ));
 sg13g2_nand2b_1 _3353_ (.Y(_1083_),
    .B(_1082_),
    .A_N(_1081_));
 sg13g2_xnor2_1 _3354_ (.Y(_1084_),
    .A(_1080_),
    .B(_1083_));
 sg13g2_nand2b_1 _3355_ (.Y(_1085_),
    .B(_1084_),
    .A_N(_1076_));
 sg13g2_nand2b_1 _3356_ (.Y(_1086_),
    .B(_1076_),
    .A_N(_1084_));
 sg13g2_and2_1 _3357_ (.A(_1085_),
    .B(_1086_),
    .X(_1087_));
 sg13g2_inv_2 _3358_ (.Y(_1088_),
    .A(_1087_));
 sg13g2_nand2_1 _3359_ (.Y(_1089_),
    .A(\videogen.fancy_shader.video_y[8] ),
    .B(net610));
 sg13g2_and2_1 _3360_ (.A(\videogen.fancy_shader.video_y[7] ),
    .B(\videogen.fancy_shader.n646[7] ),
    .X(_1090_));
 sg13g2_or2_1 _3361_ (.X(_1091_),
    .B(\videogen.fancy_shader.n646[7] ),
    .A(\videogen.fancy_shader.video_y[7] ));
 sg13g2_nand2b_1 _3362_ (.Y(_1092_),
    .B(_1091_),
    .A_N(_1090_));
 sg13g2_nor2_1 _3363_ (.A(_1083_),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_a221oi_1 _3364_ (.B2(_1080_),
    .C1(_1090_),
    .B1(_1093_),
    .A1(_1081_),
    .Y(_1094_),
    .A2(_1091_));
 sg13g2_nor2_1 _3365_ (.A(\videogen.fancy_shader.video_y[8] ),
    .B(net610),
    .Y(_1095_));
 sg13g2_xor2_1 _3366_ (.B(net610),
    .A(\videogen.fancy_shader.video_y[8] ),
    .X(_1096_));
 sg13g2_o21ai_1 _3367_ (.B1(_1089_),
    .Y(_1097_),
    .A1(_1094_),
    .A2(_1095_));
 sg13g2_xnor2_1 _3368_ (.Y(_1098_),
    .A(\videogen.fancy_shader.video_y[9] ),
    .B(\videogen.fancy_shader.n646[9] ));
 sg13g2_xnor2_1 _3369_ (.Y(_1099_),
    .A(_1097_),
    .B(_1098_));
 sg13g2_nand2_1 _3370_ (.Y(_1100_),
    .A(net610),
    .B(\videogen.fancy_shader.video_x[8] ));
 sg13g2_nor2_1 _3371_ (.A(\videogen.fancy_shader.n646[7] ),
    .B(net629),
    .Y(_1101_));
 sg13g2_xnor2_1 _3372_ (.Y(_1102_),
    .A(\videogen.fancy_shader.n646[7] ),
    .B(net629));
 sg13g2_nor2_1 _3373_ (.A(_1075_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_nor2_1 _3374_ (.A(_1074_),
    .B(_1101_),
    .Y(_1104_));
 sg13g2_a221oi_1 _3375_ (.B2(_1103_),
    .C1(_1104_),
    .B1(_1073_),
    .A1(\videogen.fancy_shader.n646[7] ),
    .Y(_1105_),
    .A2(net629));
 sg13g2_nor2_1 _3376_ (.A(net610),
    .B(\videogen.fancy_shader.video_x[8] ),
    .Y(_1106_));
 sg13g2_xor2_1 _3377_ (.B(\videogen.fancy_shader.video_x[8] ),
    .A(net610),
    .X(_1107_));
 sg13g2_o21ai_1 _3378_ (.B1(_1100_),
    .Y(_1108_),
    .A1(_1105_),
    .A2(_1106_));
 sg13g2_xor2_1 _3379_ (.B(\videogen.fancy_shader.video_x[9] ),
    .A(\videogen.fancy_shader.n646[9] ),
    .X(_1109_));
 sg13g2_xnor2_1 _3380_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_xor2_1 _3381_ (.B(_1110_),
    .A(_1099_),
    .X(_1111_));
 sg13g2_xnor2_1 _3382_ (.Y(_1112_),
    .A(_1099_),
    .B(_1110_));
 sg13g2_nand2_1 _3383_ (.Y(_1113_),
    .A(_1088_),
    .B(net542));
 sg13g2_inv_1 _3384_ (.Y(_1114_),
    .A(_1113_));
 sg13g2_nor2_1 _3385_ (.A(_1088_),
    .B(net542),
    .Y(_1115_));
 sg13g2_a21oi_1 _3386_ (.A1(_1080_),
    .A2(_1082_),
    .Y(_1116_),
    .B1(_1081_));
 sg13g2_xor2_1 _3387_ (.B(_1116_),
    .A(_1092_),
    .X(_1117_));
 sg13g2_o21ai_1 _3388_ (.B1(_1074_),
    .Y(_1118_),
    .A1(_1072_),
    .A2(_1075_));
 sg13g2_xnor2_1 _3389_ (.Y(_1119_),
    .A(_1102_),
    .B(_1118_));
 sg13g2_xnor2_1 _3390_ (.Y(_1120_),
    .A(_1117_),
    .B(_1119_));
 sg13g2_inv_1 _3391_ (.Y(_1121_),
    .A(_1120_));
 sg13g2_xnor2_1 _3392_ (.Y(_1122_),
    .A(_1105_),
    .B(_1107_));
 sg13g2_xnor2_1 _3393_ (.Y(_1123_),
    .A(_1094_),
    .B(_1096_));
 sg13g2_xnor2_1 _3394_ (.Y(_1124_),
    .A(_1122_),
    .B(_1123_));
 sg13g2_nand2_1 _3395_ (.Y(_1125_),
    .A(_1120_),
    .B(_1124_));
 sg13g2_nand3_1 _3396_ (.B(_1112_),
    .C(_1125_),
    .A(_1087_),
    .Y(_1126_));
 sg13g2_and2_1 _3397_ (.A(_1113_),
    .B(_1126_),
    .X(_1127_));
 sg13g2_nand4_1 _3398_ (.B(_1113_),
    .C(_1120_),
    .A(_1066_),
    .Y(_1128_),
    .D(_1126_));
 sg13g2_nor2_1 _3399_ (.A(_1120_),
    .B(_1124_),
    .Y(_1129_));
 sg13g2_a21oi_1 _3400_ (.A1(_1115_),
    .A2(_1120_),
    .Y(_1130_),
    .B1(_1124_));
 sg13g2_nor3_1 _3401_ (.A(_1088_),
    .B(net542),
    .C(_1125_),
    .Y(_1131_));
 sg13g2_a21oi_1 _3402_ (.A1(_1128_),
    .A2(_1130_),
    .Y(_1132_),
    .B1(_1131_));
 sg13g2_nor2_1 _3403_ (.A(_1067_),
    .B(_1132_),
    .Y(_1133_));
 sg13g2_xnor2_1 _3404_ (.Y(_1134_),
    .A(_1067_),
    .B(_1132_));
 sg13g2_nand2_1 _3405_ (.Y(_1135_),
    .A(net544),
    .B(_1127_));
 sg13g2_or2_1 _3406_ (.X(_1136_),
    .B(_1135_),
    .A(_1134_));
 sg13g2_nor3_1 _3407_ (.A(_1067_),
    .B(_1114_),
    .C(_1132_),
    .Y(_1137_));
 sg13g2_nand3b_1 _3408_ (.B(_1120_),
    .C(_1126_),
    .Y(_1138_),
    .A_N(_1137_));
 sg13g2_o21ai_1 _3409_ (.B1(_1121_),
    .Y(_1139_),
    .A1(_1115_),
    .A2(_1137_));
 sg13g2_and2_1 _3410_ (.A(_1138_),
    .B(_1139_),
    .X(_1140_));
 sg13g2_nand3_1 _3411_ (.B(_1138_),
    .C(_1139_),
    .A(_1136_),
    .Y(_1141_));
 sg13g2_a21oi_1 _3412_ (.A1(_1128_),
    .A2(_1131_),
    .Y(_1142_),
    .B1(_1130_));
 sg13g2_a21o_1 _3413_ (.A2(_1130_),
    .A1(_1128_),
    .B1(_1142_),
    .X(_1143_));
 sg13g2_inv_1 _3414_ (.Y(_1144_),
    .A(_1143_));
 sg13g2_a21oi_1 _3415_ (.A1(_1141_),
    .A2(_1143_),
    .Y(_1145_),
    .B1(_1056_));
 sg13g2_nor3_1 _3416_ (.A(net544),
    .B(_1140_),
    .C(_1144_),
    .Y(_1146_));
 sg13g2_or2_1 _3417_ (.X(_1147_),
    .B(_1146_),
    .A(_1145_));
 sg13g2_nor4_1 _3418_ (.A(_1036_),
    .B(_1134_),
    .C(_1145_),
    .D(_1146_),
    .Y(_1148_));
 sg13g2_a221oi_1 _3419_ (.B2(_1143_),
    .C1(_1134_),
    .B1(_1141_),
    .A1(_1053_),
    .Y(_1149_),
    .A2(_1054_));
 sg13g2_or3_1 _3420_ (.A(_1127_),
    .B(_1133_),
    .C(_1149_),
    .X(_1150_));
 sg13g2_o21ai_1 _3421_ (.B1(_1127_),
    .Y(_1151_),
    .A1(_1133_),
    .A2(_1149_));
 sg13g2_nand2_1 _3422_ (.Y(_1152_),
    .A(_1150_),
    .B(_1151_));
 sg13g2_a21o_2 _3423_ (.A2(_1151_),
    .A1(_1150_),
    .B1(_1148_),
    .X(_1153_));
 sg13g2_a21oi_1 _3424_ (.A1(_1136_),
    .A2(_1144_),
    .Y(_1154_),
    .B1(_1140_));
 sg13g2_a21o_2 _3425_ (.A2(_1140_),
    .A1(_1136_),
    .B1(_1154_),
    .X(_1155_));
 sg13g2_a21oi_1 _3426_ (.A1(_1153_),
    .A2(_1155_),
    .Y(_1156_),
    .B1(_1036_));
 sg13g2_nand3_1 _3427_ (.B(_1153_),
    .C(_1155_),
    .A(_1036_),
    .Y(_1157_));
 sg13g2_nand2b_1 _3428_ (.Y(_1158_),
    .B(_1157_),
    .A_N(_1156_));
 sg13g2_nor2_1 _3429_ (.A(net545),
    .B(_1147_),
    .Y(_1159_));
 sg13g2_nand3b_1 _3430_ (.B(_1157_),
    .C(_1159_),
    .Y(_1160_),
    .A_N(_1156_));
 sg13g2_a221oi_1 _3431_ (.B2(_1155_),
    .C1(_1147_),
    .B1(_1153_),
    .A1(_1032_),
    .Y(_1161_),
    .A2(_1033_));
 sg13g2_o21ai_1 _3432_ (.B1(_1134_),
    .Y(_1162_),
    .A1(_1145_),
    .A2(_1161_));
 sg13g2_or3_1 _3433_ (.A(_1134_),
    .B(_1145_),
    .C(_1161_),
    .X(_1163_));
 sg13g2_nand2_1 _3434_ (.Y(_1164_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_and3_1 _3435_ (.X(_1165_),
    .A(_1160_),
    .B(_1162_),
    .C(_1163_));
 sg13g2_nand3_1 _3436_ (.B(_1162_),
    .C(_1163_),
    .A(_1160_),
    .Y(_1166_));
 sg13g2_nor2_1 _3437_ (.A(_1148_),
    .B(_1155_),
    .Y(_1167_));
 sg13g2_o21ai_1 _3438_ (.B1(_1153_),
    .Y(_1168_),
    .A1(_1152_),
    .A2(_1167_));
 sg13g2_inv_1 _3439_ (.Y(_1169_),
    .A(_1168_));
 sg13g2_nor2_1 _3440_ (.A(_1165_),
    .B(_1169_),
    .Y(_1170_));
 sg13g2_nand3_1 _3441_ (.B(_1166_),
    .C(_1168_),
    .A(net545),
    .Y(_1171_));
 sg13g2_o21ai_1 _3442_ (.B1(_1022_),
    .Y(_1172_),
    .A1(_1165_),
    .A2(_1169_));
 sg13g2_nand2_1 _3443_ (.Y(_1173_),
    .A(_1171_),
    .B(_1172_));
 sg13g2_xnor2_1 _3444_ (.Y(_1174_),
    .A(_1004_),
    .B(_1006_));
 sg13g2_xor2_1 _3445_ (.B(_1013_),
    .A(_1012_),
    .X(_1175_));
 sg13g2_xor2_1 _3446_ (.B(_1175_),
    .A(_1174_),
    .X(_1176_));
 sg13g2_xnor2_1 _3447_ (.Y(_1177_),
    .A(_1174_),
    .B(_1175_));
 sg13g2_nand2_1 _3448_ (.Y(_1178_),
    .A(_1160_),
    .B(_1169_));
 sg13g2_a21o_1 _3449_ (.A2(_1178_),
    .A1(_1164_),
    .B1(_1165_),
    .X(_1179_));
 sg13g2_nor2_1 _3450_ (.A(_1173_),
    .B(net547),
    .Y(_1180_));
 sg13g2_nor2_1 _3451_ (.A(_1158_),
    .B(net547),
    .Y(_1181_));
 sg13g2_nand3_1 _3452_ (.B(_1172_),
    .C(_1181_),
    .A(_1171_),
    .Y(_1182_));
 sg13g2_a221oi_1 _3453_ (.B2(_1168_),
    .C1(_1158_),
    .B1(_1166_),
    .A1(_1019_),
    .Y(_1183_),
    .A2(_1020_));
 sg13g2_or3_1 _3454_ (.A(_1147_),
    .B(_1156_),
    .C(_1183_),
    .X(_1184_));
 sg13g2_o21ai_1 _3455_ (.B1(_1147_),
    .Y(_1185_),
    .A1(_1156_),
    .A2(_1183_));
 sg13g2_nand3_1 _3456_ (.B(_1184_),
    .C(_1185_),
    .A(_1182_),
    .Y(_1186_));
 sg13g2_and2_1 _3457_ (.A(_1179_),
    .B(_1186_),
    .X(_1187_));
 sg13g2_o21ai_1 _3458_ (.B1(_1173_),
    .Y(_1188_),
    .A1(net547),
    .A2(_1187_));
 sg13g2_nand3_1 _3459_ (.B(_1184_),
    .C(_1185_),
    .A(_1180_),
    .Y(_1189_));
 sg13g2_nand3_1 _3460_ (.B(net542),
    .C(_1129_),
    .A(_1088_),
    .Y(_1190_));
 sg13g2_or2_1 _3461_ (.X(_1191_),
    .B(_1129_),
    .A(net542));
 sg13g2_a21oi_1 _3462_ (.A1(_1190_),
    .A2(_1191_),
    .Y(_1192_),
    .B1(_1087_));
 sg13g2_and2_1 _3463_ (.A(_1087_),
    .B(_1191_),
    .X(_1193_));
 sg13g2_or2_1 _3464_ (.X(_1194_),
    .B(_1193_),
    .A(_1192_));
 sg13g2_inv_1 _3465_ (.Y(_1195_),
    .A(_1194_));
 sg13g2_o21ai_1 _3466_ (.B1(_1121_),
    .Y(_1196_),
    .A1(net542),
    .A2(_1124_));
 sg13g2_or4_1 _3467_ (.A(_1066_),
    .B(_1192_),
    .C(_1193_),
    .D(_1196_),
    .X(_1197_));
 sg13g2_a21oi_1 _3468_ (.A1(_1112_),
    .A2(_1121_),
    .Y(_1198_),
    .B1(_1124_));
 sg13g2_a221oi_1 _3469_ (.B2(_1191_),
    .C1(_1196_),
    .B1(_1190_),
    .A1(_1085_),
    .Y(_1199_),
    .A2(_1086_));
 sg13g2_o21ai_1 _3470_ (.B1(_1190_),
    .Y(_1200_),
    .A1(_1198_),
    .A2(_1199_));
 sg13g2_a21o_1 _3471_ (.A2(_1200_),
    .A1(_1197_),
    .B1(_1066_),
    .X(_1201_));
 sg13g2_nand2_1 _3472_ (.Y(_1202_),
    .A(_1066_),
    .B(_1200_));
 sg13g2_nand2_1 _3473_ (.Y(_1203_),
    .A(_1201_),
    .B(_1202_));
 sg13g2_inv_1 _3474_ (.Y(_1204_),
    .A(_1203_));
 sg13g2_a221oi_1 _3475_ (.B2(_1200_),
    .C1(_1194_),
    .B1(_1197_),
    .A1(_1064_),
    .Y(_1205_),
    .A2(_1065_));
 sg13g2_xnor2_1 _3476_ (.Y(_1206_),
    .A(_1195_),
    .B(_1201_));
 sg13g2_nand4_1 _3477_ (.B(_1195_),
    .C(_1201_),
    .A(_1056_),
    .Y(_1207_),
    .D(_1202_));
 sg13g2_xnor2_1 _3478_ (.Y(_1208_),
    .A(_1192_),
    .B(_1196_));
 sg13g2_o21ai_1 _3479_ (.B1(_1197_),
    .Y(_1209_),
    .A1(_1205_),
    .A2(_1208_));
 sg13g2_nor3_1 _3480_ (.A(net544),
    .B(_1203_),
    .C(_1209_),
    .Y(_1210_));
 sg13g2_o21ai_1 _3481_ (.B1(_1207_),
    .Y(_1211_),
    .A1(_1206_),
    .A2(_1210_));
 sg13g2_a21o_1 _3482_ (.A2(_1209_),
    .A1(_1207_),
    .B1(net544),
    .X(_1212_));
 sg13g2_a21oi_1 _3483_ (.A1(_1207_),
    .A2(_1209_),
    .Y(_1213_),
    .B1(net544));
 sg13g2_nand2_1 _3484_ (.Y(_1214_),
    .A(net544),
    .B(_1209_));
 sg13g2_nand2_1 _3485_ (.Y(_1215_),
    .A(_1212_),
    .B(_1214_));
 sg13g2_nand4_1 _3486_ (.B(_1204_),
    .C(_1212_),
    .A(_1036_),
    .Y(_1216_),
    .D(_1214_));
 sg13g2_a21oi_1 _3487_ (.A1(_1211_),
    .A2(_1216_),
    .Y(_1217_),
    .B1(_1037_));
 sg13g2_and2_1 _3488_ (.A(_1037_),
    .B(_1211_),
    .X(_1218_));
 sg13g2_or2_1 _3489_ (.X(_1219_),
    .B(_1218_),
    .A(_1217_));
 sg13g2_inv_1 _3490_ (.Y(_1220_),
    .A(_1219_));
 sg13g2_nor4_1 _3491_ (.A(_1022_),
    .B(_1215_),
    .C(_1217_),
    .D(_1218_),
    .Y(_1221_));
 sg13g2_a221oi_1 _3492_ (.B2(_1216_),
    .C1(_1215_),
    .B1(_1211_),
    .A1(_1034_),
    .Y(_1222_),
    .A2(_1035_));
 sg13g2_o21ai_1 _3493_ (.B1(_1203_),
    .Y(_1223_),
    .A1(_1213_),
    .A2(_1222_));
 sg13g2_nand3b_1 _3494_ (.B(_1212_),
    .C(_1204_),
    .Y(_1224_),
    .A_N(_1222_));
 sg13g2_nand3b_1 _3495_ (.B(_1223_),
    .C(_1224_),
    .Y(_1225_),
    .A_N(_1221_));
 sg13g2_nand2_1 _3496_ (.Y(_1226_),
    .A(net545),
    .B(_1225_));
 sg13g2_xnor2_1 _3497_ (.Y(_1227_),
    .A(net545),
    .B(_1225_));
 sg13g2_nor2_1 _3498_ (.A(_1219_),
    .B(_1227_),
    .Y(_1228_));
 sg13g2_xor2_1 _3499_ (.B(_1217_),
    .A(_1215_),
    .X(_1229_));
 sg13g2_nand3_1 _3500_ (.B(_1220_),
    .C(_1225_),
    .A(net545),
    .Y(_1230_));
 sg13g2_a21oi_1 _3501_ (.A1(_1229_),
    .A2(_1230_),
    .Y(_1231_),
    .B1(_1221_));
 sg13g2_o21ai_1 _3502_ (.B1(net547),
    .Y(_1232_),
    .A1(_1228_),
    .A2(_1231_));
 sg13g2_o21ai_1 _3503_ (.B1(_1226_),
    .Y(_1233_),
    .A1(_1227_),
    .A2(_1232_));
 sg13g2_xnor2_1 _3504_ (.Y(_1234_),
    .A(net609),
    .B(net630));
 sg13g2_xor2_1 _3505_ (.B(net630),
    .A(\videogen.fancy_shader.video_y[0] ),
    .X(_1235_));
 sg13g2_xnor2_1 _3506_ (.Y(_1236_),
    .A(_1219_),
    .B(_1233_));
 sg13g2_or2_1 _3507_ (.X(_1237_),
    .B(_1231_),
    .A(_1176_));
 sg13g2_nand2b_1 _3508_ (.Y(_1238_),
    .B(_1232_),
    .A_N(_1227_));
 sg13g2_a21oi_1 _3509_ (.A1(_1235_),
    .A2(_1237_),
    .Y(_1239_),
    .B1(_1238_));
 sg13g2_a221oi_1 _3510_ (.B2(_1227_),
    .C1(_1239_),
    .B1(_1237_),
    .A1(_1235_),
    .Y(_1240_),
    .A2(_1236_));
 sg13g2_nand4_1 _3511_ (.B(_1188_),
    .C(_1189_),
    .A(_1179_),
    .Y(_1241_),
    .D(_1240_));
 sg13g2_a221oi_1 _3512_ (.B2(_1186_),
    .C1(net547),
    .B1(_1179_),
    .A1(net545),
    .Y(_1242_),
    .A2(_1170_));
 sg13g2_nand2_1 _3513_ (.Y(_1243_),
    .A(_1158_),
    .B(_1172_));
 sg13g2_or2_1 _3514_ (.X(_1244_),
    .B(_1182_),
    .A(_1179_));
 sg13g2_nor2b_1 _3515_ (.A(_1183_),
    .B_N(_1244_),
    .Y(_1245_));
 sg13g2_o21ai_1 _3516_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_1242_),
    .A2(_1243_));
 sg13g2_xnor2_1 _3517_ (.Y(_1247_),
    .A(net547),
    .B(_1187_));
 sg13g2_nand3_1 _3518_ (.B(_1246_),
    .C(_1247_),
    .A(_1234_),
    .Y(_1248_));
 sg13g2_a21o_1 _3519_ (.A2(_1246_),
    .A1(_1234_),
    .B1(_1247_),
    .X(_1249_));
 sg13g2_a21o_2 _3520_ (.A2(_1249_),
    .A1(_1248_),
    .B1(_1241_),
    .X(_1250_));
 sg13g2_and2_1 _3521_ (.A(net797),
    .B(net1),
    .X(_1251_));
 sg13g2_o21ai_1 _3522_ (.B1(net619),
    .Y(_1252_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .A2(net583));
 sg13g2_nand2b_1 _3523_ (.Y(_1253_),
    .B(net624),
    .A_N(net626));
 sg13g2_nor2_1 _3524_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .B(net560),
    .Y(_1254_));
 sg13g2_nand2b_1 _3525_ (.Y(_1255_),
    .B(net627),
    .A_N(net625));
 sg13g2_nor2_1 _3526_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .B(net549),
    .Y(_1256_));
 sg13g2_nor2_1 _3527_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .B(net573),
    .Y(_1257_));
 sg13g2_nor4_1 _3528_ (.A(_1252_),
    .B(_1254_),
    .C(_1256_),
    .D(_1257_),
    .Y(_1258_));
 sg13g2_o21ai_1 _3529_ (.B1(net594),
    .Y(_1259_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .A2(net577));
 sg13g2_nor2_1 _3530_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .B(net587),
    .Y(_1260_));
 sg13g2_nor2_1 _3531_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .B(net563),
    .Y(_1261_));
 sg13g2_nor2_1 _3532_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .B(net554),
    .Y(_1262_));
 sg13g2_nor4_1 _3533_ (.A(_1259_),
    .B(_1260_),
    .C(_1261_),
    .D(_1262_),
    .Y(_1263_));
 sg13g2_nor3_1 _3534_ (.A(net616),
    .B(_1258_),
    .C(_1263_),
    .Y(_1264_));
 sg13g2_o21ai_1 _3535_ (.B1(net594),
    .Y(_1265_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .A2(net586));
 sg13g2_nor2_1 _3536_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .B(net577),
    .Y(_1266_));
 sg13g2_nor2_1 _3537_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .B(net564),
    .Y(_1267_));
 sg13g2_nor2_1 _3538_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .B(net553),
    .Y(_1268_));
 sg13g2_nor4_1 _3539_ (.A(_1265_),
    .B(_1266_),
    .C(_1267_),
    .D(_1268_),
    .Y(_1269_));
 sg13g2_o21ai_1 _3540_ (.B1(net619),
    .Y(_1270_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .A2(net572));
 sg13g2_nor2_1 _3541_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .B(net549),
    .Y(_1271_));
 sg13g2_nor2_1 _3542_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .B(net559),
    .Y(_1272_));
 sg13g2_nor2_1 _3543_ (.A(_1271_),
    .B(_1272_),
    .Y(_1273_));
 sg13g2_o21ai_1 _3544_ (.B1(_1273_),
    .Y(_1274_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ),
    .A2(net582));
 sg13g2_o21ai_1 _3545_ (.B1(net614),
    .Y(_1275_),
    .A1(_1270_),
    .A2(_1274_));
 sg13g2_o21ai_1 _3546_ (.B1(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .Y(_1276_),
    .A1(_1269_),
    .A2(_1275_));
 sg13g2_o21ai_1 _3547_ (.B1(net594),
    .Y(_1277_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .A2(net586));
 sg13g2_nor2_1 _3548_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .B(net563),
    .Y(_1278_));
 sg13g2_nor2_1 _3549_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .B(net553),
    .Y(_1279_));
 sg13g2_nor2_1 _3550_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .B(net577),
    .Y(_1280_));
 sg13g2_nor4_1 _3551_ (.A(_1277_),
    .B(_1278_),
    .C(_1279_),
    .D(_1280_),
    .Y(_1281_));
 sg13g2_o21ai_1 _3552_ (.B1(net621),
    .Y(_1282_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .A2(net578));
 sg13g2_nor2_1 _3553_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .B(net553),
    .Y(_1283_));
 sg13g2_nor2_1 _3554_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .B(net563),
    .Y(_1284_));
 sg13g2_nor2_1 _3555_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .B(net587),
    .Y(_1285_));
 sg13g2_nor4_1 _3556_ (.A(_1282_),
    .B(_1283_),
    .C(_1284_),
    .D(_1285_),
    .Y(_1286_));
 sg13g2_nor3_1 _3557_ (.A(net597),
    .B(_1281_),
    .C(_1286_),
    .Y(_1287_));
 sg13g2_nor2_1 _3558_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .B(net589),
    .Y(_1288_));
 sg13g2_nor2_1 _3559_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .B(net566),
    .Y(_1289_));
 sg13g2_nor2_1 _3560_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .B(net556),
    .Y(_1290_));
 sg13g2_o21ai_1 _3561_ (.B1(net622),
    .Y(_1291_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .A2(net580));
 sg13g2_nor4_1 _3562_ (.A(_1288_),
    .B(_1289_),
    .C(_1290_),
    .D(_1291_),
    .Y(_1292_));
 sg13g2_o21ai_1 _3563_ (.B1(net594),
    .Y(_1293_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .A2(net566));
 sg13g2_nor2_1 _3564_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .B(net589),
    .Y(_1294_));
 sg13g2_nor2_1 _3565_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .B(net556),
    .Y(_1295_));
 sg13g2_nor2_1 _3566_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .B(net580),
    .Y(_1296_));
 sg13g2_nor4_1 _3567_ (.A(_1293_),
    .B(_1294_),
    .C(_1295_),
    .D(_1296_),
    .Y(_1297_));
 sg13g2_nor3_1 _3568_ (.A(net618),
    .B(_1292_),
    .C(_1297_),
    .Y(_1298_));
 sg13g2_nor3_1 _3569_ (.A(net613),
    .B(_1287_),
    .C(_1298_),
    .Y(_1299_));
 sg13g2_nor2_1 _3570_ (.A(_0636_),
    .B(_1299_),
    .Y(_1300_));
 sg13g2_o21ai_1 _3571_ (.B1(_1300_),
    .Y(_1301_),
    .A1(_1264_),
    .A2(_1276_));
 sg13g2_o21ai_1 _3572_ (.B1(net622),
    .Y(_1302_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .A2(net588));
 sg13g2_nor2_1 _3573_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .B(net565),
    .Y(_1303_));
 sg13g2_nor2_1 _3574_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .B(net555),
    .Y(_1304_));
 sg13g2_nor2_1 _3575_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .B(net579),
    .Y(_1305_));
 sg13g2_nor4_1 _3576_ (.A(_1302_),
    .B(_1303_),
    .C(_1304_),
    .D(_1305_),
    .Y(_1306_));
 sg13g2_nor2_1 _3577_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .B(net579),
    .Y(_1307_));
 sg13g2_nor2_1 _3578_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .B(net555),
    .Y(_1308_));
 sg13g2_nor2_1 _3579_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .B(net588),
    .Y(_1309_));
 sg13g2_o21ai_1 _3580_ (.B1(net594),
    .Y(_1310_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .A2(net565));
 sg13g2_nor4_1 _3581_ (.A(_1307_),
    .B(_1308_),
    .C(_1309_),
    .D(_1310_),
    .Y(_1311_));
 sg13g2_nor3_1 _3582_ (.A(net618),
    .B(_1306_),
    .C(_1311_),
    .Y(_1312_));
 sg13g2_o21ai_1 _3583_ (.B1(net593),
    .Y(_1313_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .A2(net562));
 sg13g2_nor2_1 _3584_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .B(net585),
    .Y(_1314_));
 sg13g2_nor2_1 _3585_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .B(net575),
    .Y(_1315_));
 sg13g2_nor2_1 _3586_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .B(net551),
    .Y(_1316_));
 sg13g2_nor4_1 _3587_ (.A(_1313_),
    .B(_1314_),
    .C(_1315_),
    .D(_1316_),
    .Y(_1317_));
 sg13g2_o21ai_1 _3588_ (.B1(net620),
    .Y(_1318_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .A2(net585));
 sg13g2_nor2_1 _3589_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .B(net574),
    .Y(_1319_));
 sg13g2_nor2_1 _3590_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .B(net561),
    .Y(_1320_));
 sg13g2_nor2_1 _3591_ (.A(_1319_),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_o21ai_1 _3592_ (.B1(_1321_),
    .Y(_1322_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .A2(net551));
 sg13g2_o21ai_1 _3593_ (.B1(net615),
    .Y(_1323_),
    .A1(_1318_),
    .A2(_1322_));
 sg13g2_o21ai_1 _3594_ (.B1(net612),
    .Y(_1324_),
    .A1(_1317_),
    .A2(_1323_));
 sg13g2_o21ai_1 _3595_ (.B1(net593),
    .Y(_1325_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .A2(net561));
 sg13g2_nor2_1 _3596_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .B(net574),
    .Y(_1326_));
 sg13g2_nor2_1 _3597_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .B(net584),
    .Y(_1327_));
 sg13g2_nor2_1 _3598_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .B(net552),
    .Y(_1328_));
 sg13g2_nor4_1 _3599_ (.A(_1325_),
    .B(_1326_),
    .C(_1327_),
    .D(_1328_),
    .Y(_1329_));
 sg13g2_o21ai_1 _3600_ (.B1(net619),
    .Y(_1330_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .A2(net582));
 sg13g2_nor2_1 _3601_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .B(net549),
    .Y(_1331_));
 sg13g2_nor2_1 _3602_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .B(net559),
    .Y(_1332_));
 sg13g2_nor2_1 _3603_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .B(net572),
    .Y(_1333_));
 sg13g2_nor4_1 _3604_ (.A(_1330_),
    .B(_1331_),
    .C(_1332_),
    .D(_1333_),
    .Y(_1334_));
 sg13g2_nor3_1 _3605_ (.A(net599),
    .B(_1329_),
    .C(_1334_),
    .Y(_1335_));
 sg13g2_o21ai_1 _3606_ (.B1(net623),
    .Y(_1336_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .A2(net562));
 sg13g2_nor2_1 _3607_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .B(net585),
    .Y(_1337_));
 sg13g2_nor2_1 _3608_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .B(net551),
    .Y(_1338_));
 sg13g2_nor2_1 _3609_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .B(net575),
    .Y(_1339_));
 sg13g2_nor4_1 _3610_ (.A(_1336_),
    .B(_1337_),
    .C(_1338_),
    .D(_1339_),
    .Y(_1340_));
 sg13g2_o21ai_1 _3611_ (.B1(net593),
    .Y(_1341_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .A2(net574));
 sg13g2_nor2_1 _3612_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .B(net552),
    .Y(_1342_));
 sg13g2_nor2_1 _3613_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .B(net561),
    .Y(_1343_));
 sg13g2_nor2_1 _3614_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .B(net584),
    .Y(_1344_));
 sg13g2_nor4_1 _3615_ (.A(_1341_),
    .B(_1342_),
    .C(_1343_),
    .D(_1344_),
    .Y(_1345_));
 sg13g2_nor3_1 _3616_ (.A(net614),
    .B(_1340_),
    .C(_1345_),
    .Y(_1346_));
 sg13g2_nor3_1 _3617_ (.A(net612),
    .B(_1335_),
    .C(_1346_),
    .Y(_1347_));
 sg13g2_nor2_1 _3618_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_o21ai_1 _3619_ (.B1(_1348_),
    .Y(_1349_),
    .A1(_1312_),
    .A2(_1324_));
 sg13g2_nand3_1 _3620_ (.B(_1301_),
    .C(_1349_),
    .A(net2),
    .Y(_1350_));
 sg13g2_o21ai_1 _3621_ (.B1(_1350_),
    .Y(_1351_),
    .A1(net2),
    .A2(_0651_));
 sg13g2_inv_4 _3622_ (.A(_1351_),
    .Y(_1352_));
 sg13g2_o21ai_1 _3623_ (.B1(net618),
    .Y(_1353_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ),
    .A2(net575));
 sg13g2_nor2_1 _3624_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .B(net555),
    .Y(_1354_));
 sg13g2_nor2_1 _3625_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .B(net588),
    .Y(_1355_));
 sg13g2_nor2_1 _3626_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .B(net565),
    .Y(_1356_));
 sg13g2_nor4_1 _3627_ (.A(_1353_),
    .B(_1354_),
    .C(_1355_),
    .D(_1356_),
    .Y(_1357_));
 sg13g2_o21ai_1 _3628_ (.B1(net598),
    .Y(_1358_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .A2(net555));
 sg13g2_nor2_1 _3629_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .B(net579),
    .Y(_1359_));
 sg13g2_nor2_1 _3630_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ),
    .B(net588),
    .Y(_1360_));
 sg13g2_nor2_1 _3631_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .B(net565),
    .Y(_1361_));
 sg13g2_nor4_1 _3632_ (.A(_1358_),
    .B(_1359_),
    .C(_1360_),
    .D(_1361_),
    .Y(_1362_));
 sg13g2_nor3_1 _3633_ (.A(net622),
    .B(_1357_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_o21ai_1 _3634_ (.B1(net615),
    .Y(_1364_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .A2(net562));
 sg13g2_nor2_1 _3635_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .B(net585),
    .Y(_1365_));
 sg13g2_nor2_1 _3636_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .B(net575),
    .Y(_1366_));
 sg13g2_nor2_1 _3637_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .B(net551),
    .Y(_1367_));
 sg13g2_nor4_1 _3638_ (.A(_1364_),
    .B(_1365_),
    .C(_1366_),
    .D(_1367_),
    .Y(_1368_));
 sg13g2_o21ai_1 _3639_ (.B1(net596),
    .Y(_1369_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .A2(net562));
 sg13g2_nor2_1 _3640_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .B(net584),
    .Y(_1370_));
 sg13g2_nor2_1 _3641_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .B(net551),
    .Y(_1371_));
 sg13g2_nor2_1 _3642_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .B(net575),
    .Y(_1372_));
 sg13g2_nor4_1 _3643_ (.A(_1369_),
    .B(_1370_),
    .C(_1371_),
    .D(_1372_),
    .Y(_1373_));
 sg13g2_nor3_1 _3644_ (.A(net592),
    .B(_1368_),
    .C(_1373_),
    .Y(_1374_));
 sg13g2_nand2b_1 _3645_ (.Y(_1375_),
    .B(net613),
    .A_N(_1374_));
 sg13g2_o21ai_1 _3646_ (.B1(net614),
    .Y(_1376_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .A2(net582));
 sg13g2_nor2_1 _3647_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .B(net549),
    .Y(_1377_));
 sg13g2_nor2_1 _3648_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .B(net559),
    .Y(_1378_));
 sg13g2_nor2_1 _3649_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .B(net572),
    .Y(_1379_));
 sg13g2_nor4_1 _3650_ (.A(_1376_),
    .B(_1377_),
    .C(_1378_),
    .D(_1379_),
    .Y(_1380_));
 sg13g2_o21ai_1 _3651_ (.B1(net596),
    .Y(_1381_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .A2(net583));
 sg13g2_nor2_1 _3652_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .B(net559),
    .Y(_1382_));
 sg13g2_nor2_1 _3653_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .B(net573),
    .Y(_1383_));
 sg13g2_nor2_1 _3654_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .B(net550),
    .Y(_1384_));
 sg13g2_nor4_1 _3655_ (.A(_1381_),
    .B(_1382_),
    .C(_1383_),
    .D(_1384_),
    .Y(_1385_));
 sg13g2_nor3_1 _3656_ (.A(net592),
    .B(_1380_),
    .C(_1385_),
    .Y(_1386_));
 sg13g2_o21ai_1 _3657_ (.B1(net615),
    .Y(_1387_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .A2(net552));
 sg13g2_nor2_1 _3658_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ),
    .B(net574),
    .Y(_1388_));
 sg13g2_nor2_1 _3659_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .B(net584),
    .Y(_1389_));
 sg13g2_nor2_1 _3660_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .B(net561),
    .Y(_1390_));
 sg13g2_nor4_1 _3661_ (.A(_1387_),
    .B(_1388_),
    .C(_1389_),
    .D(_1390_),
    .Y(_1391_));
 sg13g2_o21ai_1 _3662_ (.B1(net596),
    .Y(_1392_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .A2(net574));
 sg13g2_nor2_1 _3663_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .B(net561),
    .Y(_1393_));
 sg13g2_nor2_1 _3664_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .B(net552),
    .Y(_1394_));
 sg13g2_nor2_1 _3665_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ),
    .B(net584),
    .Y(_1395_));
 sg13g2_nor4_1 _3666_ (.A(_1392_),
    .B(_1393_),
    .C(_1394_),
    .D(_1395_),
    .Y(_1396_));
 sg13g2_nor3_1 _3667_ (.A(net620),
    .B(_1391_),
    .C(_1396_),
    .Y(_1397_));
 sg13g2_nor3_1 _3668_ (.A(net612),
    .B(_1386_),
    .C(_1397_),
    .Y(_1398_));
 sg13g2_nor2_1 _3669_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_o21ai_1 _3670_ (.B1(_1399_),
    .Y(_1400_),
    .A1(_1363_),
    .A2(_1375_));
 sg13g2_o21ai_1 _3671_ (.B1(net597),
    .Y(_1401_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .A2(net563));
 sg13g2_nor2_1 _3672_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ),
    .B(net578),
    .Y(_1402_));
 sg13g2_nor2_1 _3673_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .B(net554),
    .Y(_1403_));
 sg13g2_nor2_1 _3674_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .B(net587),
    .Y(_1404_));
 sg13g2_nor4_1 _3675_ (.A(_1401_),
    .B(_1402_),
    .C(_1403_),
    .D(_1404_),
    .Y(_1405_));
 sg13g2_o21ai_1 _3676_ (.B1(net617),
    .Y(_1406_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .A2(net586));
 sg13g2_nor2_1 _3677_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .B(net577),
    .Y(_1407_));
 sg13g2_nor2_1 _3678_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .B(net564),
    .Y(_1408_));
 sg13g2_nor2_1 _3679_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ),
    .B(net553),
    .Y(_1409_));
 sg13g2_nor4_1 _3680_ (.A(_1406_),
    .B(_1407_),
    .C(_1408_),
    .D(_1409_),
    .Y(_1410_));
 sg13g2_nor3_1 _3681_ (.A(net621),
    .B(_1405_),
    .C(_1410_),
    .Y(_1411_));
 sg13g2_o21ai_1 _3682_ (.B1(net614),
    .Y(_1412_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ),
    .A2(net572));
 sg13g2_nor2_1 _3683_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .B(net549),
    .Y(_1413_));
 sg13g2_nor2_1 _3684_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .B(net559),
    .Y(_1414_));
 sg13g2_nor2_1 _3685_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ),
    .B(net582),
    .Y(_1415_));
 sg13g2_nor4_1 _3686_ (.A(_1412_),
    .B(_1413_),
    .C(_1414_),
    .D(_1415_),
    .Y(_1416_));
 sg13g2_o21ai_1 _3687_ (.B1(net596),
    .Y(_1417_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .A2(net560));
 sg13g2_nor2_1 _3688_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .B(net573),
    .Y(_1418_));
 sg13g2_nor2_1 _3689_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .B(net550),
    .Y(_1419_));
 sg13g2_nor2_1 _3690_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .B(net583),
    .Y(_1420_));
 sg13g2_nor4_1 _3691_ (.A(_1417_),
    .B(_1418_),
    .C(_1419_),
    .D(_1420_),
    .Y(_1421_));
 sg13g2_nor3_1 _3692_ (.A(net592),
    .B(_1416_),
    .C(_1421_),
    .Y(_1422_));
 sg13g2_nor3_1 _3693_ (.A(_0637_),
    .B(_1411_),
    .C(_1422_),
    .Y(_1423_));
 sg13g2_o21ai_1 _3694_ (.B1(net597),
    .Y(_1424_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .A2(net590));
 sg13g2_nor2_1 _3695_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .B(net556),
    .Y(_1425_));
 sg13g2_nor2_1 _3696_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .B(net566),
    .Y(_1426_));
 sg13g2_nor2_1 _3697_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .B(net579),
    .Y(_1427_));
 sg13g2_nor4_1 _3698_ (.A(_1424_),
    .B(_1425_),
    .C(_1426_),
    .D(_1427_),
    .Y(_1428_));
 sg13g2_o21ai_1 _3699_ (.B1(net616),
    .Y(_1429_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .A2(net578));
 sg13g2_nor2_1 _3700_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .B(net563),
    .Y(_1430_));
 sg13g2_nor2_1 _3701_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .B(net553),
    .Y(_1431_));
 sg13g2_nor2_1 _3702_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .B(net586),
    .Y(_1432_));
 sg13g2_nor4_1 _3703_ (.A(_1429_),
    .B(_1430_),
    .C(_1431_),
    .D(_1432_),
    .Y(_1433_));
 sg13g2_nor3_1 _3704_ (.A(net594),
    .B(_1428_),
    .C(_1433_),
    .Y(_1434_));
 sg13g2_o21ai_1 _3705_ (.B1(net618),
    .Y(_1435_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .A2(net577));
 sg13g2_nor2_1 _3706_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .B(net565),
    .Y(_1436_));
 sg13g2_nor2_1 _3707_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .B(net586),
    .Y(_1437_));
 sg13g2_nor2_1 _3708_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ),
    .B(net553),
    .Y(_1438_));
 sg13g2_nor4_1 _3709_ (.A(_1435_),
    .B(_1436_),
    .C(_1437_),
    .D(_1438_),
    .Y(_1439_));
 sg13g2_o21ai_1 _3710_ (.B1(net597),
    .Y(_1440_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .A2(net567));
 sg13g2_nor2_1 _3711_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .B(net589),
    .Y(_1441_));
 sg13g2_nor2_1 _3712_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .B(net556),
    .Y(_1442_));
 sg13g2_nor2_1 _3713_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ),
    .B(net580),
    .Y(_1443_));
 sg13g2_nor4_1 _3714_ (.A(_1440_),
    .B(_1441_),
    .C(_1442_),
    .D(_1443_),
    .Y(_1444_));
 sg13g2_nor3_1 _3715_ (.A(net622),
    .B(_1439_),
    .C(_1444_),
    .Y(_1445_));
 sg13g2_nor3_1 _3716_ (.A(net613),
    .B(_1434_),
    .C(_1445_),
    .Y(_1446_));
 sg13g2_nor3_1 _3717_ (.A(_0636_),
    .B(_1423_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_nor2_1 _3718_ (.A(_0650_),
    .B(_1447_),
    .Y(_1448_));
 sg13g2_a22oi_1 _3719_ (.Y(_1449_),
    .B1(_1400_),
    .B2(_1448_),
    .A2(_0650_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[1] ));
 sg13g2_nand2_1 _3720_ (.Y(_1450_),
    .A(_1352_),
    .B(_1449_));
 sg13g2_nor2_1 _3721_ (.A(net749),
    .B(net1),
    .Y(_1451_));
 sg13g2_o21ai_1 _3722_ (.B1(net618),
    .Y(_1452_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .A2(net565));
 sg13g2_nor2_1 _3723_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .B(net555),
    .Y(_1453_));
 sg13g2_nor2_1 _3724_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ),
    .B(net579),
    .Y(_1454_));
 sg13g2_nor2_1 _3725_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .B(net588),
    .Y(_1455_));
 sg13g2_nor4_1 _3726_ (.A(_1452_),
    .B(_1453_),
    .C(_1454_),
    .D(_1455_),
    .Y(_1456_));
 sg13g2_o21ai_1 _3727_ (.B1(net598),
    .Y(_1457_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .A2(net555));
 sg13g2_nor2_1 _3728_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .B(net579),
    .Y(_1458_));
 sg13g2_nor2_1 _3729_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .B(net565),
    .Y(_1459_));
 sg13g2_nor2_1 _3730_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ),
    .B(net589),
    .Y(_1460_));
 sg13g2_nor4_1 _3731_ (.A(_1457_),
    .B(_1458_),
    .C(_1459_),
    .D(_1460_),
    .Y(_1461_));
 sg13g2_nor3_1 _3732_ (.A(net622),
    .B(_1456_),
    .C(_1461_),
    .Y(_1462_));
 sg13g2_o21ai_1 _3733_ (.B1(net596),
    .Y(_1463_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .A2(net562));
 sg13g2_nor2_1 _3734_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .B(net551),
    .Y(_1464_));
 sg13g2_nor2_1 _3735_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .B(net584),
    .Y(_1465_));
 sg13g2_nor2_1 _3736_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .B(net575),
    .Y(_1466_));
 sg13g2_nor4_1 _3737_ (.A(_1463_),
    .B(_1464_),
    .C(_1465_),
    .D(_1466_),
    .Y(_1467_));
 sg13g2_o21ai_1 _3738_ (.B1(net615),
    .Y(_1468_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .A2(net551));
 sg13g2_nor2_1 _3739_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .B(net574),
    .Y(_1469_));
 sg13g2_nor2_1 _3740_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .B(net561),
    .Y(_1470_));
 sg13g2_nor2_1 _3741_ (.A(_1469_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_o21ai_1 _3742_ (.B1(_1471_),
    .Y(_1472_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .A2(net585));
 sg13g2_o21ai_1 _3743_ (.B1(net620),
    .Y(_1473_),
    .A1(_1468_),
    .A2(_1472_));
 sg13g2_o21ai_1 _3744_ (.B1(net613),
    .Y(_1474_),
    .A1(_1467_),
    .A2(_1473_));
 sg13g2_o21ai_1 _3745_ (.B1(net596),
    .Y(_1475_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .A2(net572));
 sg13g2_nor2_1 _3746_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .B(net559),
    .Y(_1476_));
 sg13g2_nor2_1 _3747_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .B(net549),
    .Y(_1477_));
 sg13g2_nor2_1 _3748_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .B(net582),
    .Y(_1478_));
 sg13g2_nor4_1 _3749_ (.A(_1475_),
    .B(_1476_),
    .C(_1477_),
    .D(_1478_),
    .Y(_1479_));
 sg13g2_o21ai_1 _3750_ (.B1(net614),
    .Y(_1480_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .A2(net549));
 sg13g2_nor2_1 _3751_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .B(net572),
    .Y(_1481_));
 sg13g2_nor2_1 _3752_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .B(net559),
    .Y(_1482_));
 sg13g2_nor2_1 _3753_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .B(net582),
    .Y(_1483_));
 sg13g2_nor4_1 _3754_ (.A(_1480_),
    .B(_1481_),
    .C(_1482_),
    .D(_1483_),
    .Y(_1484_));
 sg13g2_nor3_1 _3755_ (.A(net592),
    .B(_1479_),
    .C(_1484_),
    .Y(_1485_));
 sg13g2_o21ai_1 _3756_ (.B1(net615),
    .Y(_1486_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .A2(net561));
 sg13g2_nor2_1 _3757_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ),
    .B(net584),
    .Y(_1487_));
 sg13g2_nor2_1 _3758_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .B(net574),
    .Y(_1488_));
 sg13g2_nor2_1 _3759_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .B(net552),
    .Y(_1489_));
 sg13g2_nor4_1 _3760_ (.A(_1486_),
    .B(_1487_),
    .C(_1488_),
    .D(_1489_),
    .Y(_1490_));
 sg13g2_o21ai_1 _3761_ (.B1(net599),
    .Y(_1491_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .A2(net552));
 sg13g2_nor2_1 _3762_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ),
    .B(net574),
    .Y(_1492_));
 sg13g2_nor2_1 _3763_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .B(net562),
    .Y(_1493_));
 sg13g2_nor2_1 _3764_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .B(net584),
    .Y(_1494_));
 sg13g2_nor4_1 _3765_ (.A(_1491_),
    .B(_1492_),
    .C(_1493_),
    .D(_1494_),
    .Y(_1495_));
 sg13g2_nor3_1 _3766_ (.A(net620),
    .B(_1490_),
    .C(_1495_),
    .Y(_1496_));
 sg13g2_nor3_1 _3767_ (.A(net612),
    .B(_1485_),
    .C(_1496_),
    .Y(_1497_));
 sg13g2_nor2_1 _3768_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_o21ai_1 _3769_ (.B1(_1498_),
    .Y(_1499_),
    .A1(_1462_),
    .A2(_1474_));
 sg13g2_o21ai_1 _3770_ (.B1(net617),
    .Y(_1500_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .A2(net586));
 sg13g2_nor2_1 _3771_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .B(net577),
    .Y(_1501_));
 sg13g2_nor2_1 _3772_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .B(net564),
    .Y(_1502_));
 sg13g2_nor2_1 _3773_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .B(net553),
    .Y(_1503_));
 sg13g2_nor4_1 _3774_ (.A(_1500_),
    .B(_1501_),
    .C(_1502_),
    .D(_1503_),
    .Y(_1504_));
 sg13g2_o21ai_1 _3775_ (.B1(net597),
    .Y(_1505_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .A2(net554));
 sg13g2_nor2_1 _3776_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .B(net563),
    .Y(_1506_));
 sg13g2_nor2_1 _3777_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .B(net587),
    .Y(_1507_));
 sg13g2_nor2_1 _3778_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .B(net581),
    .Y(_1508_));
 sg13g2_nor4_1 _3779_ (.A(_1505_),
    .B(_1506_),
    .C(_1507_),
    .D(_1508_),
    .Y(_1509_));
 sg13g2_nor3_1 _3780_ (.A(net621),
    .B(_1504_),
    .C(_1509_),
    .Y(_1510_));
 sg13g2_o21ai_1 _3781_ (.B1(net614),
    .Y(_1511_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ),
    .A2(net572));
 sg13g2_nor2_1 _3782_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .B(net559),
    .Y(_1512_));
 sg13g2_nor2_1 _3783_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .B(net582),
    .Y(_1513_));
 sg13g2_nor2_1 _3784_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .B(net549),
    .Y(_1514_));
 sg13g2_nor4_1 _3785_ (.A(_1511_),
    .B(_1512_),
    .C(_1513_),
    .D(_1514_),
    .Y(_1515_));
 sg13g2_o21ai_1 _3786_ (.B1(net596),
    .Y(_1516_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .A2(net583));
 sg13g2_nor2_1 _3787_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .B(net573),
    .Y(_1517_));
 sg13g2_nor2_1 _3788_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .B(net560),
    .Y(_1518_));
 sg13g2_nor2_1 _3789_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .B(net550),
    .Y(_1519_));
 sg13g2_nor4_1 _3790_ (.A(_1516_),
    .B(_1517_),
    .C(_1518_),
    .D(_1519_),
    .Y(_1520_));
 sg13g2_nor3_1 _3791_ (.A(net592),
    .B(_1515_),
    .C(_1520_),
    .Y(_1521_));
 sg13g2_nor3_1 _3792_ (.A(_0637_),
    .B(_1510_),
    .C(_1521_),
    .Y(_1522_));
 sg13g2_o21ai_1 _3793_ (.B1(net597),
    .Y(_1523_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .A2(net566));
 sg13g2_nor2_1 _3794_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .B(net580),
    .Y(_1524_));
 sg13g2_nor2_1 _3795_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .B(net589),
    .Y(_1525_));
 sg13g2_nor2_1 _3796_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .B(net556),
    .Y(_1526_));
 sg13g2_nor4_1 _3797_ (.A(_1523_),
    .B(_1524_),
    .C(_1525_),
    .D(_1526_),
    .Y(_1527_));
 sg13g2_o21ai_1 _3798_ (.B1(net616),
    .Y(_1528_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ),
    .A2(net578));
 sg13g2_nor2_1 _3799_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ),
    .B(net586),
    .Y(_1529_));
 sg13g2_nor2_1 _3800_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .B(net563),
    .Y(_1530_));
 sg13g2_nor2_1 _3801_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .B(net554),
    .Y(_1531_));
 sg13g2_nor4_1 _3802_ (.A(_1528_),
    .B(_1529_),
    .C(_1530_),
    .D(_1531_),
    .Y(_1532_));
 sg13g2_nor3_1 _3803_ (.A(net594),
    .B(_1527_),
    .C(_1532_),
    .Y(_1533_));
 sg13g2_o21ai_1 _3804_ (.B1(net617),
    .Y(_1534_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .A2(net577));
 sg13g2_nor2_1 _3805_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .B(net554),
    .Y(_1535_));
 sg13g2_nor2_1 _3806_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .B(net586),
    .Y(_1536_));
 sg13g2_nor2_1 _3807_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .B(net564),
    .Y(_1537_));
 sg13g2_nor4_1 _3808_ (.A(_1534_),
    .B(_1535_),
    .C(_1536_),
    .D(_1537_),
    .Y(_1538_));
 sg13g2_o21ai_1 _3809_ (.B1(net598),
    .Y(_1539_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .A2(net556));
 sg13g2_nor2_1 _3810_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .B(net580),
    .Y(_1540_));
 sg13g2_nor2_1 _3811_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .B(net589),
    .Y(_1541_));
 sg13g2_nor2_1 _3812_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .B(net566),
    .Y(_1542_));
 sg13g2_nor4_1 _3813_ (.A(_1539_),
    .B(_1540_),
    .C(_1541_),
    .D(_1542_),
    .Y(_1543_));
 sg13g2_nor3_1 _3814_ (.A(net622),
    .B(_1538_),
    .C(_1543_),
    .Y(_1544_));
 sg13g2_nor3_1 _3815_ (.A(net613),
    .B(_1533_),
    .C(_1544_),
    .Y(_1545_));
 sg13g2_nor3_1 _3816_ (.A(_0636_),
    .B(_1522_),
    .C(_1545_),
    .Y(_1546_));
 sg13g2_nor2_1 _3817_ (.A(_0650_),
    .B(_1546_),
    .Y(_1547_));
 sg13g2_a22oi_1 _3818_ (.Y(_1548_),
    .B1(_1499_),
    .B2(_1547_),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A1(_0650_));
 sg13g2_nor2b_2 _3819_ (.A(_1548_),
    .B_N(_1451_),
    .Y(_1549_));
 sg13g2_inv_1 _3820_ (.Y(_1550_),
    .A(_1549_));
 sg13g2_a22oi_1 _3821_ (.Y(_1551_),
    .B1(_1450_),
    .B2(_1549_),
    .A2(_1251_),
    .A1(_1250_));
 sg13g2_inv_1 _3822_ (.Y(_0372_),
    .A(_1551_));
 sg13g2_nor2_1 _3823_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .B(net565),
    .Y(_1552_));
 sg13g2_nor2_1 _3824_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .B(net579),
    .Y(_1553_));
 sg13g2_nor2_1 _3825_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .B(net555),
    .Y(_1554_));
 sg13g2_o21ai_1 _3826_ (.B1(net620),
    .Y(_1555_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .A2(net588));
 sg13g2_nor4_1 _3827_ (.A(_1552_),
    .B(_1553_),
    .C(_1554_),
    .D(_1555_),
    .Y(_1556_));
 sg13g2_nor2_1 _3828_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .B(net555),
    .Y(_1557_));
 sg13g2_nor2_1 _3829_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ),
    .B(net588),
    .Y(_1558_));
 sg13g2_nor2_1 _3830_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .B(net566),
    .Y(_1559_));
 sg13g2_o21ai_1 _3831_ (.B1(net595),
    .Y(_1560_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .A2(net579));
 sg13g2_nor4_1 _3832_ (.A(_1557_),
    .B(_1558_),
    .C(_1559_),
    .D(_1560_),
    .Y(_1561_));
 sg13g2_or2_1 _3833_ (.X(_1562_),
    .B(net562),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ));
 sg13g2_nand2b_1 _3834_ (.Y(_1563_),
    .B(_0674_),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ));
 sg13g2_or2_1 _3835_ (.X(_1564_),
    .B(net575),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ));
 sg13g2_or2_1 _3836_ (.X(_1565_),
    .B(net561),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ));
 sg13g2_or2_1 _3837_ (.X(_1566_),
    .B(net573),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ));
 sg13g2_nand2b_1 _3838_ (.Y(_1567_),
    .B(_0674_),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ));
 sg13g2_o21ai_1 _3839_ (.B1(_1567_),
    .Y(_1568_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .A2(net560));
 sg13g2_or2_1 _3840_ (.X(_1569_),
    .B(net553),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ));
 sg13g2_or2_1 _3841_ (.X(_1570_),
    .B(net563),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ));
 sg13g2_o21ai_1 _3842_ (.B1(net622),
    .Y(_1571_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .A2(net580));
 sg13g2_nor2_1 _3843_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .B(net556),
    .Y(_1572_));
 sg13g2_nor2_1 _3844_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .B(net566),
    .Y(_1573_));
 sg13g2_nor2_1 _3845_ (.A(_1572_),
    .B(_1573_),
    .Y(_1574_));
 sg13g2_o21ai_1 _3846_ (.B1(_1574_),
    .Y(_1575_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .A2(net589));
 sg13g2_nor2_1 _3847_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .B(net590),
    .Y(_1576_));
 sg13g2_nor2_1 _3848_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .B(net556),
    .Y(_1577_));
 sg13g2_o21ai_1 _3849_ (.B1(net595),
    .Y(_1578_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .A2(net567));
 sg13g2_nor3_1 _3850_ (.A(_1576_),
    .B(_1577_),
    .C(_1578_),
    .Y(_1579_));
 sg13g2_o21ai_1 _3851_ (.B1(_1579_),
    .Y(_1580_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ),
    .A2(net580));
 sg13g2_or2_1 _3852_ (.X(_1581_),
    .B(net2),
    .A(\videogen.test_lut_thingy.gol_counter_reg[0] ));
 sg13g2_mux4_1 _3853_ (.S0(net627),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .S1(net624),
    .X(_1582_));
 sg13g2_mux4_1 _3854_ (.S0(net626),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .S1(net625),
    .X(_1583_));
 sg13g2_mux2_1 _3855_ (.A0(_1582_),
    .A1(_1583_),
    .S(net594),
    .X(_1584_));
 sg13g2_o21ai_1 _3856_ (.B1(_1566_),
    .Y(_1585_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .A2(net550));
 sg13g2_o21ai_1 _3857_ (.B1(net620),
    .Y(_1586_),
    .A1(_1568_),
    .A2(_1585_));
 sg13g2_mux4_1 _3858_ (.S0(net625),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .S1(net628),
    .X(_1587_));
 sg13g2_o21ai_1 _3859_ (.B1(_1586_),
    .Y(_1588_),
    .A1(net621),
    .A2(_1587_));
 sg13g2_o21ai_1 _3860_ (.B1(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .Y(_1589_),
    .A1(net616),
    .A2(_1588_));
 sg13g2_a21oi_1 _3861_ (.A1(net616),
    .A2(_1584_),
    .Y(_1590_),
    .B1(_1589_));
 sg13g2_o21ai_1 _3862_ (.B1(_1569_),
    .Y(_1591_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .A2(net578));
 sg13g2_o21ai_1 _3863_ (.B1(_1570_),
    .Y(_1592_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .A2(net587));
 sg13g2_o21ai_1 _3864_ (.B1(net621),
    .Y(_1593_),
    .A1(_1591_),
    .A2(_1592_));
 sg13g2_mux4_1 _3865_ (.S0(net625),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .S1(net628),
    .X(_1594_));
 sg13g2_nor2_1 _3866_ (.A(net621),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_nor2_1 _3867_ (.A(net597),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_o21ai_1 _3868_ (.B1(_1580_),
    .Y(_1597_),
    .A1(_1571_),
    .A2(_1575_));
 sg13g2_a221oi_1 _3869_ (.B2(net597),
    .C1(net613),
    .B1(_1597_),
    .A1(_1593_),
    .Y(_1598_),
    .A2(_1596_));
 sg13g2_nor3_1 _3870_ (.A(_0636_),
    .B(_1590_),
    .C(_1598_),
    .Y(_1599_));
 sg13g2_mux4_1 _3871_ (.S0(net624),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .S1(net627),
    .X(_1600_));
 sg13g2_mux4_1 _3872_ (.S0(net627),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .S1(net624),
    .X(_1601_));
 sg13g2_mux4_1 _3873_ (.S0(net627),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .S1(net624),
    .X(_1602_));
 sg13g2_mux4_1 _3874_ (.S0(net624),
    .A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .A2(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .A3(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .S1(net627),
    .X(_1603_));
 sg13g2_mux4_1 _3875_ (.S0(net623),
    .A0(_1600_),
    .A1(_1601_),
    .A2(_1603_),
    .A3(_1602_),
    .S1(net599),
    .X(_1604_));
 sg13g2_o21ai_1 _3876_ (.B1(_1563_),
    .Y(_1605_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .A2(net573));
 sg13g2_o21ai_1 _3877_ (.B1(_1562_),
    .Y(_1606_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .A2(net551));
 sg13g2_o21ai_1 _3878_ (.B1(net593),
    .Y(_1607_),
    .A1(_1605_),
    .A2(_1606_));
 sg13g2_o21ai_1 _3879_ (.B1(_1565_),
    .Y(_1608_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .A2(net552));
 sg13g2_o21ai_1 _3880_ (.B1(_1564_),
    .Y(_1609_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .A2(net585));
 sg13g2_o21ai_1 _3881_ (.B1(net620),
    .Y(_1610_),
    .A1(_1608_),
    .A2(_1609_));
 sg13g2_nand3_1 _3882_ (.B(_1607_),
    .C(_1610_),
    .A(net615),
    .Y(_1611_));
 sg13g2_o21ai_1 _3883_ (.B1(net598),
    .Y(_1612_),
    .A1(_1556_),
    .A2(_1561_));
 sg13g2_nand3_1 _3884_ (.B(_1611_),
    .C(_1612_),
    .A(net612),
    .Y(_1613_));
 sg13g2_o21ai_1 _3885_ (.B1(_1613_),
    .Y(_1614_),
    .A1(net612),
    .A2(_1604_));
 sg13g2_o21ai_1 _3886_ (.B1(net2),
    .Y(_1615_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .A2(_1614_));
 sg13g2_o21ai_1 _3887_ (.B1(_1581_),
    .Y(_1616_),
    .A1(_1599_),
    .A2(_1615_));
 sg13g2_nand2b_1 _3888_ (.Y(_1617_),
    .B(_1616_),
    .A_N(_1449_));
 sg13g2_a21oi_1 _3889_ (.A1(net1),
    .A2(_1250_),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_nor2_1 _3890_ (.A(_1551_),
    .B(_1618_),
    .Y(_0374_));
 sg13g2_a21oi_1 _3891_ (.A1(_1351_),
    .A2(_1618_),
    .Y(_0373_),
    .B1(_1551_));
 sg13g2_nand2_1 _3892_ (.Y(_1619_),
    .A(_1449_),
    .B(_1616_));
 sg13g2_nand3_1 _3893_ (.B(_1449_),
    .C(_1616_),
    .A(_1352_),
    .Y(_1620_));
 sg13g2_and2_1 _3894_ (.A(_1549_),
    .B(_1620_),
    .X(_1621_));
 sg13g2_a21o_1 _3895_ (.A2(_1251_),
    .A1(_1250_),
    .B1(_1621_),
    .X(_0375_));
 sg13g2_xor2_1 _3896_ (.B(\videogen.fancy_shader.n646[0] ),
    .A(\videogen.fancy_shader.video_y[0] ),
    .X(_1622_));
 sg13g2_nand2_2 _3897_ (.Y(_1623_),
    .A(_1006_),
    .B(_1622_));
 sg13g2_o21ai_1 _3898_ (.B1(_1623_),
    .Y(_1624_),
    .A1(_1174_),
    .A2(_1622_));
 sg13g2_xnor2_1 _3899_ (.Y(_1625_),
    .A(_1175_),
    .B(_1624_));
 sg13g2_nor2_2 _3900_ (.A(_1010_),
    .B(_1623_),
    .Y(_1626_));
 sg13g2_nand2_1 _3901_ (.Y(_1627_),
    .A(_1036_),
    .B(_1626_));
 sg13g2_or2_1 _3902_ (.X(_1628_),
    .B(_1626_),
    .A(_1036_));
 sg13g2_and2_1 _3903_ (.A(_1627_),
    .B(_1628_),
    .X(_1629_));
 sg13g2_nand2_1 _3904_ (.Y(_1630_),
    .A(net546),
    .B(_1626_));
 sg13g2_nand3_1 _3905_ (.B(_1052_),
    .C(_1626_),
    .A(net546),
    .Y(_1631_));
 sg13g2_and4_1 _3906_ (.A(net546),
    .B(_1052_),
    .C(_1063_),
    .D(_1626_),
    .X(_1632_));
 sg13g2_xnor2_1 _3907_ (.Y(_1633_),
    .A(_1063_),
    .B(_1631_));
 sg13g2_xor2_1 _3908_ (.B(_1633_),
    .A(_1060_),
    .X(_1634_));
 sg13g2_inv_2 _3909_ (.Y(_1635_),
    .A(_1634_));
 sg13g2_and2_1 _3910_ (.A(_1093_),
    .B(_1632_),
    .X(_1636_));
 sg13g2_xnor2_1 _3911_ (.Y(_1637_),
    .A(_1124_),
    .B(_1636_));
 sg13g2_nand2_1 _3912_ (.Y(_1638_),
    .A(_1123_),
    .B(_1636_));
 sg13g2_xnor2_1 _3913_ (.Y(_1639_),
    .A(_1112_),
    .B(_1638_));
 sg13g2_xnor2_1 _3914_ (.Y(_1640_),
    .A(net542),
    .B(_1638_));
 sg13g2_xnor2_1 _3915_ (.Y(_1641_),
    .A(_1087_),
    .B(_1632_));
 sg13g2_nand2_1 _3916_ (.Y(_1642_),
    .A(_1084_),
    .B(_1632_));
 sg13g2_xor2_1 _3917_ (.B(_1642_),
    .A(_1120_),
    .X(_1643_));
 sg13g2_or3_1 _3918_ (.A(_1640_),
    .B(_1641_),
    .C(_1643_),
    .X(_1644_));
 sg13g2_and2_1 _3919_ (.A(_1637_),
    .B(_1644_),
    .X(_1645_));
 sg13g2_nor3_1 _3920_ (.A(_1637_),
    .B(_1641_),
    .C(_1643_),
    .Y(_1646_));
 sg13g2_nor3_2 _3921_ (.A(_1640_),
    .B(_1641_),
    .C(_1646_),
    .Y(_1647_));
 sg13g2_xor2_1 _3922_ (.B(_1647_),
    .A(_1643_),
    .X(_1648_));
 sg13g2_and2_1 _3923_ (.A(_1640_),
    .B(_1641_),
    .X(_1649_));
 sg13g2_nor2_1 _3924_ (.A(_1647_),
    .B(_1649_),
    .Y(_1650_));
 sg13g2_inv_1 _3925_ (.Y(_1651_),
    .A(_1650_));
 sg13g2_nand2_1 _3926_ (.Y(_1652_),
    .A(_1634_),
    .B(_1650_));
 sg13g2_nor4_1 _3927_ (.A(_1635_),
    .B(_1643_),
    .C(_1647_),
    .D(_1649_),
    .Y(_1653_));
 sg13g2_or4_1 _3928_ (.A(_1635_),
    .B(_1643_),
    .C(_1647_),
    .D(_1649_),
    .X(_1654_));
 sg13g2_nor2_1 _3929_ (.A(_1637_),
    .B(_1644_),
    .Y(_1655_));
 sg13g2_a21oi_2 _3930_ (.B1(_1655_),
    .Y(_1656_),
    .A2(_1654_),
    .A1(_1645_));
 sg13g2_xnor2_1 _3931_ (.Y(_1657_),
    .A(_1634_),
    .B(_1656_));
 sg13g2_xnor2_1 _3932_ (.Y(_1658_),
    .A(_1635_),
    .B(_1656_));
 sg13g2_xor2_1 _3933_ (.B(_1630_),
    .A(net544),
    .X(_1659_));
 sg13g2_inv_1 _3934_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_nor2_1 _3935_ (.A(_1651_),
    .B(_1659_),
    .Y(_1661_));
 sg13g2_nand2_1 _3936_ (.Y(_1662_),
    .A(_1657_),
    .B(_1661_));
 sg13g2_o21ai_1 _3937_ (.B1(_1648_),
    .Y(_1663_),
    .A1(_1652_),
    .A2(_1656_));
 sg13g2_nand2_1 _3938_ (.Y(_1664_),
    .A(_1653_),
    .B(_1655_));
 sg13g2_nand2_1 _3939_ (.Y(_1665_),
    .A(_1663_),
    .B(_1664_));
 sg13g2_a22oi_1 _3940_ (.Y(_1666_),
    .B1(_1663_),
    .B2(_1664_),
    .A2(_1661_),
    .A1(_1657_));
 sg13g2_nor2_1 _3941_ (.A(_1653_),
    .B(_1655_),
    .Y(_1667_));
 sg13g2_nor2_1 _3942_ (.A(_1645_),
    .B(_1654_),
    .Y(_1668_));
 sg13g2_nor2_1 _3943_ (.A(_1667_),
    .B(_1668_),
    .Y(_1669_));
 sg13g2_a21oi_1 _3944_ (.A1(_1662_),
    .A2(_1669_),
    .Y(_1670_),
    .B1(_1665_));
 sg13g2_or2_1 _3945_ (.X(_1671_),
    .B(_1670_),
    .A(_1666_));
 sg13g2_o21ai_1 _3946_ (.B1(_1660_),
    .Y(_1672_),
    .A1(_1666_),
    .A2(_1669_));
 sg13g2_inv_1 _3947_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_or3_1 _3948_ (.A(_1660_),
    .B(_1666_),
    .C(_1669_),
    .X(_1674_));
 sg13g2_nand2_1 _3949_ (.Y(_1675_),
    .A(_1672_),
    .B(_1674_));
 sg13g2_nor2_1 _3950_ (.A(_1629_),
    .B(_1658_),
    .Y(_1676_));
 sg13g2_and3_1 _3951_ (.X(_1677_),
    .A(_1672_),
    .B(_1674_),
    .C(_1676_));
 sg13g2_o21ai_1 _3952_ (.B1(_1651_),
    .Y(_1678_),
    .A1(_1635_),
    .A2(_1656_));
 sg13g2_o21ai_1 _3953_ (.B1(_1678_),
    .Y(_1679_),
    .A1(_1652_),
    .A2(_1656_));
 sg13g2_o21ai_1 _3954_ (.B1(_1679_),
    .Y(_1680_),
    .A1(_1658_),
    .A2(_1672_));
 sg13g2_or3_1 _3955_ (.A(_1658_),
    .B(_1672_),
    .C(_1679_),
    .X(_1681_));
 sg13g2_and2_1 _3956_ (.A(_1680_),
    .B(_1681_),
    .X(_1682_));
 sg13g2_a21o_1 _3957_ (.A2(_1681_),
    .A1(_1680_),
    .B1(_1677_),
    .X(_1683_));
 sg13g2_a21o_1 _3958_ (.A2(_1683_),
    .A1(_1671_),
    .B1(_1629_),
    .X(_1684_));
 sg13g2_nand3_1 _3959_ (.B(_1671_),
    .C(_1682_),
    .A(_1629_),
    .Y(_1685_));
 sg13g2_and2_1 _3960_ (.A(_1684_),
    .B(_1685_),
    .X(_1686_));
 sg13g2_xnor2_1 _3961_ (.Y(_1687_),
    .A(net545),
    .B(_1623_));
 sg13g2_xor2_1 _3962_ (.B(_1623_),
    .A(_1021_),
    .X(_1688_));
 sg13g2_nor2_1 _3963_ (.A(_1675_),
    .B(_1687_),
    .Y(_1689_));
 sg13g2_nand3_1 _3964_ (.B(_1685_),
    .C(_1689_),
    .A(_1684_),
    .Y(_1690_));
 sg13g2_a221oi_1 _3965_ (.B2(_1683_),
    .C1(_1675_),
    .B1(_1671_),
    .A1(_1627_),
    .Y(_1691_),
    .A2(_1628_));
 sg13g2_nand3b_1 _3966_ (.B(_1657_),
    .C(_1672_),
    .Y(_1692_),
    .A_N(_1691_));
 sg13g2_o21ai_1 _3967_ (.B1(_1658_),
    .Y(_1693_),
    .A1(_1673_),
    .A2(_1691_));
 sg13g2_nand2_1 _3968_ (.Y(_1694_),
    .A(_1692_),
    .B(_1693_));
 sg13g2_nand3_1 _3969_ (.B(_1692_),
    .C(_1693_),
    .A(_1690_),
    .Y(_1695_));
 sg13g2_o21ai_1 _3970_ (.B1(_1682_),
    .Y(_1696_),
    .A1(_1671_),
    .A2(_1677_));
 sg13g2_nand2_1 _3971_ (.Y(_1697_),
    .A(_1683_),
    .B(_1696_));
 sg13g2_a21oi_1 _3972_ (.A1(_1695_),
    .A2(_1697_),
    .Y(_1698_),
    .B1(_1687_));
 sg13g2_nand2_1 _3973_ (.Y(_1699_),
    .A(_1686_),
    .B(_1698_));
 sg13g2_or2_1 _3974_ (.X(_1700_),
    .B(_1698_),
    .A(_1686_));
 sg13g2_a21o_1 _3975_ (.A2(_1700_),
    .A1(_1699_),
    .B1(_1234_),
    .X(_1701_));
 sg13g2_nor2_1 _3976_ (.A(_1625_),
    .B(_1701_),
    .Y(_1702_));
 sg13g2_xnor2_1 _3977_ (.Y(_1703_),
    .A(_1675_),
    .B(_1684_));
 sg13g2_xnor2_1 _3978_ (.Y(_1704_),
    .A(_1699_),
    .B(_1703_));
 sg13g2_a21oi_1 _3979_ (.A1(_1625_),
    .A2(_1701_),
    .Y(_1705_),
    .B1(_1704_));
 sg13g2_nor2b_1 _3980_ (.A(_1702_),
    .B_N(_1705_),
    .Y(_1706_));
 sg13g2_nand3_1 _3981_ (.B(_1694_),
    .C(_1697_),
    .A(_1687_),
    .Y(_1707_));
 sg13g2_nor2b_1 _3982_ (.A(_1698_),
    .B_N(_1707_),
    .Y(_1708_));
 sg13g2_nand3_1 _3983_ (.B(_1701_),
    .C(_1704_),
    .A(_1625_),
    .Y(_1709_));
 sg13g2_nand2_1 _3984_ (.Y(_1710_),
    .A(_1708_),
    .B(_1709_));
 sg13g2_mux2_1 _3985_ (.A0(_1694_),
    .A1(_1697_),
    .S(_1690_),
    .X(_1711_));
 sg13g2_a21oi_1 _3986_ (.A1(_1702_),
    .A2(_1704_),
    .Y(_1712_),
    .B1(_1708_));
 sg13g2_nand2_1 _3987_ (.Y(_1713_),
    .A(_1240_),
    .B(_1711_));
 sg13g2_nor2_1 _3988_ (.A(_1712_),
    .B(_1713_),
    .Y(_1714_));
 sg13g2_o21ai_1 _3989_ (.B1(_1714_),
    .Y(_1715_),
    .A1(_1706_),
    .A2(_1710_));
 sg13g2_nand2_1 _3990_ (.Y(_1716_),
    .A(_1251_),
    .B(_1715_));
 sg13g2_nor2_1 _3991_ (.A(_1352_),
    .B(_1548_),
    .Y(_1717_));
 sg13g2_o21ai_1 _3992_ (.B1(_1451_),
    .Y(_1718_),
    .A1(_1352_),
    .A2(_1548_));
 sg13g2_a21o_1 _3993_ (.A2(_1548_),
    .A1(_1352_),
    .B1(_1718_),
    .X(_1719_));
 sg13g2_nand2_1 _3994_ (.Y(_0377_),
    .A(_1716_),
    .B(_1719_));
 sg13g2_or2_1 _3995_ (.X(_1720_),
    .B(_1616_),
    .A(_1449_));
 sg13g2_or2_1 _3996_ (.X(_1721_),
    .B(_1720_),
    .A(_1718_));
 sg13g2_nand3_1 _3997_ (.B(_1719_),
    .C(_1721_),
    .A(_1716_),
    .Y(_0376_));
 sg13g2_and2_1 _3998_ (.A(_1619_),
    .B(_1717_),
    .X(_1722_));
 sg13g2_a21oi_1 _3999_ (.A1(_1450_),
    .A2(_1451_),
    .Y(_1723_),
    .B1(_1549_));
 sg13g2_o21ai_1 _4000_ (.B1(_1716_),
    .Y(_0378_),
    .A1(_1722_),
    .A2(_1723_));
 sg13g2_xnor2_1 _4001_ (.Y(_1724_),
    .A(\videogen.fancy_shader.n646[0] ),
    .B(\videogen.fancy_shader.video_x[0] ));
 sg13g2_or2_1 _4002_ (.X(_1725_),
    .B(_1724_),
    .A(_1013_));
 sg13g2_nor2_2 _4003_ (.A(_1039_),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_inv_1 _4004_ (.Y(_1727_),
    .A(_1726_));
 sg13g2_xnor2_1 _4005_ (.Y(_1728_),
    .A(_1659_),
    .B(_1726_));
 sg13g2_nor3_2 _4006_ (.A(_1039_),
    .B(_1068_),
    .C(_1725_),
    .Y(_1729_));
 sg13g2_nand2_1 _4007_ (.Y(_1730_),
    .A(_1076_),
    .B(_1729_));
 sg13g2_xnor2_1 _4008_ (.Y(_1731_),
    .A(_1076_),
    .B(_1729_));
 sg13g2_xnor2_1 _4009_ (.Y(_1732_),
    .A(_1084_),
    .B(_1632_));
 sg13g2_nand2b_1 _4010_ (.Y(_1733_),
    .B(_1732_),
    .A_N(_1731_));
 sg13g2_nand2b_1 _4011_ (.Y(_1734_),
    .B(_1731_),
    .A_N(_1732_));
 sg13g2_and2_1 _4012_ (.A(_1733_),
    .B(_1734_),
    .X(_1735_));
 sg13g2_xor2_1 _4013_ (.B(_1730_),
    .A(_1643_),
    .X(_1736_));
 sg13g2_and2_1 _4014_ (.A(_1103_),
    .B(_1729_),
    .X(_1737_));
 sg13g2_nand2_1 _4015_ (.Y(_1738_),
    .A(_1122_),
    .B(_1737_));
 sg13g2_xnor2_1 _4016_ (.Y(_1739_),
    .A(_1639_),
    .B(_1738_));
 sg13g2_nand2b_1 _4017_ (.Y(_1740_),
    .B(_1739_),
    .A_N(_1736_));
 sg13g2_xor2_1 _4018_ (.B(_1737_),
    .A(_1637_),
    .X(_1741_));
 sg13g2_inv_1 _4019_ (.Y(_1742_),
    .A(_1741_));
 sg13g2_a21oi_1 _4020_ (.A1(_1739_),
    .A2(_1741_),
    .Y(_1743_),
    .B1(_1736_));
 sg13g2_inv_1 _4021_ (.Y(_1744_),
    .A(_1743_));
 sg13g2_a221oi_1 _4022_ (.B2(_1741_),
    .C1(_1736_),
    .B1(_1739_),
    .A1(_1733_),
    .Y(_1745_),
    .A2(_1734_));
 sg13g2_nor4_1 _4023_ (.A(_1735_),
    .B(_1736_),
    .C(_1739_),
    .D(_1742_),
    .Y(_1746_));
 sg13g2_o21ai_1 _4024_ (.B1(_1739_),
    .Y(_1747_),
    .A1(_1736_),
    .A2(_1742_));
 sg13g2_nor2b_1 _4025_ (.A(_1746_),
    .B_N(_1747_),
    .Y(_1748_));
 sg13g2_xor2_1 _4026_ (.B(_1748_),
    .A(_1735_),
    .X(_1749_));
 sg13g2_nand2_1 _4027_ (.Y(_1750_),
    .A(_1046_),
    .B(_1726_));
 sg13g2_a21oi_1 _4028_ (.A1(_1060_),
    .A2(_1750_),
    .Y(_1751_),
    .B1(_1729_));
 sg13g2_xnor2_1 _4029_ (.Y(_1752_),
    .A(_1633_),
    .B(_1751_));
 sg13g2_nor2_1 _4030_ (.A(_1744_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_nand2_1 _4031_ (.Y(_1754_),
    .A(_1740_),
    .B(_1741_));
 sg13g2_o21ai_1 _4032_ (.B1(_1745_),
    .Y(_1755_),
    .A1(_1739_),
    .A2(_1741_));
 sg13g2_a21o_1 _4033_ (.A2(_1755_),
    .A1(_1754_),
    .B1(_1746_),
    .X(_1756_));
 sg13g2_a221oi_1 _4034_ (.B2(_1755_),
    .C1(_1752_),
    .B1(_1754_),
    .A1(_1741_),
    .Y(_1757_),
    .A2(_1745_));
 sg13g2_o21ai_1 _4035_ (.B1(_1749_),
    .Y(_1758_),
    .A1(_1753_),
    .A2(_1757_));
 sg13g2_o21ai_1 _4036_ (.B1(_1744_),
    .Y(_1759_),
    .A1(_1735_),
    .A2(_1748_));
 sg13g2_nand2_1 _4037_ (.Y(_1760_),
    .A(_1755_),
    .B(_1759_));
 sg13g2_a22oi_1 _4038_ (.Y(_1761_),
    .B1(_1758_),
    .B2(_1760_),
    .A2(_1753_),
    .A1(_1749_));
 sg13g2_a221oi_1 _4039_ (.B2(_1752_),
    .C1(_1757_),
    .B1(_1756_),
    .A1(_1749_),
    .Y(_1762_),
    .A2(_1753_));
 sg13g2_nor2b_1 _4040_ (.A(_1728_),
    .B_N(_1749_),
    .Y(_1763_));
 sg13g2_or2_1 _4041_ (.X(_1764_),
    .B(_1757_),
    .A(_1749_));
 sg13g2_and2_1 _4042_ (.A(_1762_),
    .B(_1763_),
    .X(_1765_));
 sg13g2_nor2_2 _4043_ (.A(_1761_),
    .B(_1765_),
    .Y(_1766_));
 sg13g2_nor2_1 _4044_ (.A(_1728_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_xor2_1 _4045_ (.B(_1766_),
    .A(_1728_),
    .X(_1768_));
 sg13g2_xnor2_1 _4046_ (.Y(_1769_),
    .A(_1728_),
    .B(_1766_));
 sg13g2_nor2_1 _4047_ (.A(_1018_),
    .B(_1725_),
    .Y(_1770_));
 sg13g2_o21ai_1 _4048_ (.B1(_1727_),
    .Y(_1771_),
    .A1(_1027_),
    .A2(_1770_));
 sg13g2_xor2_1 _4049_ (.B(_1626_),
    .A(net546),
    .X(_1772_));
 sg13g2_xnor2_1 _4050_ (.Y(_1773_),
    .A(_1771_),
    .B(_1772_));
 sg13g2_nand3_1 _4051_ (.B(_1768_),
    .C(_1773_),
    .A(_1762_),
    .Y(_1774_));
 sg13g2_a22oi_1 _4052_ (.Y(_1775_),
    .B1(_1767_),
    .B2(_1762_),
    .A2(_1764_),
    .A1(_1758_));
 sg13g2_o21ai_1 _4053_ (.B1(_1774_),
    .Y(_1776_),
    .A1(_1765_),
    .A2(_1775_));
 sg13g2_nand2_1 _4054_ (.Y(_1777_),
    .A(_1773_),
    .B(_1776_));
 sg13g2_xor2_1 _4055_ (.B(_1776_),
    .A(_1773_),
    .X(_1778_));
 sg13g2_xnor2_1 _4056_ (.Y(_1779_),
    .A(_1688_),
    .B(_1725_));
 sg13g2_nand2b_1 _4057_ (.Y(_1780_),
    .B(_1778_),
    .A_N(_1779_));
 sg13g2_xnor2_1 _4058_ (.Y(_1781_),
    .A(_1762_),
    .B(_1767_));
 sg13g2_nand2b_1 _4059_ (.Y(_1782_),
    .B(_1774_),
    .A_N(_1781_));
 sg13g2_or2_1 _4060_ (.X(_1783_),
    .B(_1780_),
    .A(_1769_));
 sg13g2_o21ai_1 _4061_ (.B1(_1781_),
    .Y(_1784_),
    .A1(_1769_),
    .A2(_1777_));
 sg13g2_nand2_1 _4062_ (.Y(_1785_),
    .A(_1774_),
    .B(_1784_));
 sg13g2_a21oi_1 _4063_ (.A1(_1783_),
    .A2(_1785_),
    .Y(_1786_),
    .B1(_1779_));
 sg13g2_a21oi_1 _4064_ (.A1(_1769_),
    .A2(_1782_),
    .Y(_1787_),
    .B1(_1780_));
 sg13g2_a21oi_1 _4065_ (.A1(_1773_),
    .A2(_1776_),
    .Y(_1788_),
    .B1(_1787_));
 sg13g2_xnor2_1 _4066_ (.Y(_1789_),
    .A(_1769_),
    .B(_1788_));
 sg13g2_nand2_1 _4067_ (.Y(_1790_),
    .A(_1234_),
    .B(_1778_));
 sg13g2_a21o_1 _4068_ (.A2(_1790_),
    .A1(_1789_),
    .B1(_1177_),
    .X(_1791_));
 sg13g2_a21oi_1 _4069_ (.A1(_1779_),
    .A2(_1785_),
    .Y(_1792_),
    .B1(_1786_));
 sg13g2_nor2_1 _4070_ (.A(net547),
    .B(_1234_),
    .Y(_1793_));
 sg13g2_o21ai_1 _4071_ (.B1(_1793_),
    .Y(_1794_),
    .A1(_1778_),
    .A2(_1789_));
 sg13g2_nand3_1 _4072_ (.B(_1792_),
    .C(_1794_),
    .A(_1791_),
    .Y(_1795_));
 sg13g2_xor2_1 _4073_ (.B(_1725_),
    .A(_1174_),
    .X(_1796_));
 sg13g2_nor2b_1 _4074_ (.A(_1010_),
    .B_N(_1174_),
    .Y(_1797_));
 sg13g2_xnor2_1 _4075_ (.Y(_1798_),
    .A(_1021_),
    .B(_1796_));
 sg13g2_and2_1 _4076_ (.A(_1031_),
    .B(_1797_),
    .X(_1799_));
 sg13g2_xnor2_1 _4077_ (.Y(_1800_),
    .A(_1726_),
    .B(_1799_));
 sg13g2_nand2_1 _4078_ (.Y(_1801_),
    .A(_1052_),
    .B(_1799_));
 sg13g2_xnor2_1 _4079_ (.Y(_1802_),
    .A(_1055_),
    .B(_1800_));
 sg13g2_inv_1 _4080_ (.Y(_1803_),
    .A(_1802_));
 sg13g2_nand3_1 _4081_ (.B(_1063_),
    .C(_1799_),
    .A(_1052_),
    .Y(_1804_));
 sg13g2_xor2_1 _4082_ (.B(_1801_),
    .A(_1063_),
    .X(_1805_));
 sg13g2_xnor2_1 _4083_ (.Y(_1806_),
    .A(_1751_),
    .B(_1805_));
 sg13g2_and4_1 _4084_ (.A(_1052_),
    .B(_1063_),
    .C(_1084_),
    .D(_1799_),
    .X(_1807_));
 sg13g2_nand2_1 _4085_ (.Y(_1808_),
    .A(_1117_),
    .B(_1807_));
 sg13g2_xor2_1 _4086_ (.B(_1808_),
    .A(_1737_),
    .X(_1809_));
 sg13g2_nand3_1 _4087_ (.B(_1123_),
    .C(_1807_),
    .A(_1117_),
    .Y(_1810_));
 sg13g2_xnor2_1 _4088_ (.Y(_1811_),
    .A(_1124_),
    .B(_1809_));
 sg13g2_xor2_1 _4089_ (.B(_1804_),
    .A(_1084_),
    .X(_1812_));
 sg13g2_xnor2_1 _4090_ (.Y(_1813_),
    .A(_1731_),
    .B(_1812_));
 sg13g2_xor2_1 _4091_ (.B(_1812_),
    .A(_1731_),
    .X(_1814_));
 sg13g2_xor2_1 _4092_ (.B(_1810_),
    .A(_1738_),
    .X(_1815_));
 sg13g2_nand2_1 _4093_ (.Y(_1816_),
    .A(net542),
    .B(_1815_));
 sg13g2_nand2b_1 _4094_ (.Y(_1817_),
    .B(_1112_),
    .A_N(_1815_));
 sg13g2_xnor2_1 _4095_ (.Y(_1818_),
    .A(_1111_),
    .B(_1815_));
 sg13g2_xnor2_1 _4096_ (.Y(_1819_),
    .A(_1730_),
    .B(_1807_));
 sg13g2_xor2_1 _4097_ (.B(_1819_),
    .A(_1120_),
    .X(_1820_));
 sg13g2_inv_1 _4098_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_nand3_1 _4099_ (.B(_1818_),
    .C(_1820_),
    .A(_1813_),
    .Y(_1822_));
 sg13g2_nor2b_1 _4100_ (.A(_1822_),
    .B_N(_1811_),
    .Y(_1823_));
 sg13g2_a221oi_1 _4101_ (.B2(_1811_),
    .C1(_1814_),
    .B1(_1820_),
    .A1(_1816_),
    .Y(_1824_),
    .A2(_1817_));
 sg13g2_nor2_1 _4102_ (.A(_1813_),
    .B(_1818_),
    .Y(_1825_));
 sg13g2_or2_1 _4103_ (.X(_1826_),
    .B(_1825_),
    .A(_1824_));
 sg13g2_or4_1 _4104_ (.A(_1806_),
    .B(_1821_),
    .C(_1824_),
    .D(_1825_),
    .X(_1827_));
 sg13g2_nor2b_1 _4105_ (.A(_1811_),
    .B_N(_1822_),
    .Y(_1828_));
 sg13g2_a21oi_1 _4106_ (.A1(_1827_),
    .A2(_1828_),
    .Y(_1829_),
    .B1(_1823_));
 sg13g2_xnor2_1 _4107_ (.Y(_1830_),
    .A(_1806_),
    .B(_1829_));
 sg13g2_nor2_1 _4108_ (.A(_1803_),
    .B(_1830_),
    .Y(_1831_));
 sg13g2_or3_1 _4109_ (.A(_1803_),
    .B(_1826_),
    .C(_1830_),
    .X(_1832_));
 sg13g2_nor3_1 _4110_ (.A(_1806_),
    .B(_1826_),
    .C(_1829_),
    .Y(_1833_));
 sg13g2_xnor2_1 _4111_ (.Y(_1834_),
    .A(_1821_),
    .B(_1824_));
 sg13g2_xnor2_1 _4112_ (.Y(_1835_),
    .A(_1833_),
    .B(_1834_));
 sg13g2_mux2_1 _4113_ (.A0(_1828_),
    .A1(_1823_),
    .S(_1827_),
    .X(_1836_));
 sg13g2_a21o_2 _4114_ (.A2(_1835_),
    .A1(_1832_),
    .B1(_1836_),
    .X(_1837_));
 sg13g2_nand2_1 _4115_ (.Y(_1838_),
    .A(_1802_),
    .B(_1837_));
 sg13g2_xnor2_1 _4116_ (.Y(_1839_),
    .A(_1803_),
    .B(_1837_));
 sg13g2_xnor2_1 _4117_ (.Y(_1840_),
    .A(_1802_),
    .B(_1837_));
 sg13g2_xor2_1 _4118_ (.B(_1797_),
    .A(_1031_),
    .X(_1841_));
 sg13g2_xnor2_1 _4119_ (.Y(_1842_),
    .A(_1771_),
    .B(_1841_));
 sg13g2_inv_1 _4120_ (.Y(_1843_),
    .A(_1842_));
 sg13g2_nor2_1 _4121_ (.A(_1830_),
    .B(_1842_),
    .Y(_1844_));
 sg13g2_nand2_1 _4122_ (.Y(_1845_),
    .A(_1839_),
    .B(_1844_));
 sg13g2_o21ai_1 _4123_ (.B1(_1826_),
    .Y(_1846_),
    .A1(_1806_),
    .A2(_1829_));
 sg13g2_nor2b_1 _4124_ (.A(_1833_),
    .B_N(_1846_),
    .Y(_1847_));
 sg13g2_a21o_1 _4125_ (.A2(_1837_),
    .A1(_1831_),
    .B1(_1847_),
    .X(_1848_));
 sg13g2_nand3_1 _4126_ (.B(_1837_),
    .C(_1847_),
    .A(_1831_),
    .Y(_1849_));
 sg13g2_and2_1 _4127_ (.A(_1848_),
    .B(_1849_),
    .X(_1850_));
 sg13g2_a22oi_1 _4128_ (.Y(_1851_),
    .B1(_1848_),
    .B2(_1849_),
    .A2(_1844_),
    .A1(_1839_));
 sg13g2_a21oi_1 _4129_ (.A1(_1832_),
    .A2(_1836_),
    .Y(_1852_),
    .B1(_1835_));
 sg13g2_a21oi_1 _4130_ (.A1(_1832_),
    .A2(_1835_),
    .Y(_1853_),
    .B1(_1852_));
 sg13g2_o21ai_1 _4131_ (.B1(_1843_),
    .Y(_1854_),
    .A1(_1851_),
    .A2(_1853_));
 sg13g2_nand3b_1 _4132_ (.B(_1850_),
    .C(_1842_),
    .Y(_1855_),
    .A_N(_1853_));
 sg13g2_and2_1 _4133_ (.A(_1854_),
    .B(_1855_),
    .X(_1856_));
 sg13g2_nand2_1 _4134_ (.Y(_1857_),
    .A(_1854_),
    .B(_1855_));
 sg13g2_nor2_1 _4135_ (.A(_1798_),
    .B(_1857_),
    .Y(_1858_));
 sg13g2_nor2_1 _4136_ (.A(_1798_),
    .B(_1840_),
    .Y(_1859_));
 sg13g2_and3_1 _4137_ (.X(_1860_),
    .A(_1854_),
    .B(_1855_),
    .C(_1859_));
 sg13g2_xnor2_1 _4138_ (.Y(_1861_),
    .A(_1830_),
    .B(_1838_));
 sg13g2_o21ai_1 _4139_ (.B1(_1861_),
    .Y(_1862_),
    .A1(_1840_),
    .A2(_1854_));
 sg13g2_or3_1 _4140_ (.A(_1840_),
    .B(_1854_),
    .C(_1861_),
    .X(_1863_));
 sg13g2_nand2_1 _4141_ (.Y(_1864_),
    .A(_1862_),
    .B(_1863_));
 sg13g2_a21oi_1 _4142_ (.A1(_1862_),
    .A2(_1863_),
    .Y(_1865_),
    .B1(_1860_));
 sg13g2_a21o_1 _4143_ (.A2(_1863_),
    .A1(_1862_),
    .B1(_1860_),
    .X(_1866_));
 sg13g2_o21ai_1 _4144_ (.B1(_1845_),
    .Y(_1867_),
    .A1(_1851_),
    .A2(_1853_));
 sg13g2_a21oi_1 _4145_ (.A1(_1850_),
    .A2(_1867_),
    .Y(_1868_),
    .B1(_1851_));
 sg13g2_a21o_1 _4146_ (.A2(_1867_),
    .A1(_1850_),
    .B1(_1851_),
    .X(_1869_));
 sg13g2_a21oi_1 _4147_ (.A1(_1866_),
    .A2(_1869_),
    .Y(_1870_),
    .B1(_1798_));
 sg13g2_and3_1 _4148_ (.X(_1871_),
    .A(_1798_),
    .B(_1866_),
    .C(_1869_));
 sg13g2_nor2_1 _4149_ (.A(_1870_),
    .B(_1871_),
    .Y(_1872_));
 sg13g2_nand2b_1 _4150_ (.Y(_1873_),
    .B(_1724_),
    .A_N(_1175_));
 sg13g2_nand2_1 _4151_ (.Y(_1874_),
    .A(_1725_),
    .B(_1873_));
 sg13g2_xor2_1 _4152_ (.B(_1874_),
    .A(_1174_),
    .X(_1875_));
 sg13g2_nor4_1 _4153_ (.A(_1857_),
    .B(_1870_),
    .C(_1871_),
    .D(_1875_),
    .Y(_1876_));
 sg13g2_xnor2_1 _4154_ (.Y(_1877_),
    .A(_1839_),
    .B(_1854_));
 sg13g2_o21ai_1 _4155_ (.B1(_1858_),
    .Y(_1878_),
    .A1(_1865_),
    .A2(_1868_));
 sg13g2_xnor2_1 _4156_ (.Y(_1879_),
    .A(_1877_),
    .B(_1878_));
 sg13g2_nor2_1 _4157_ (.A(_1876_),
    .B(_1879_),
    .Y(_1880_));
 sg13g2_a21oi_1 _4158_ (.A1(_1866_),
    .A2(_1869_),
    .Y(_1881_),
    .B1(_1860_));
 sg13g2_o21ai_1 _4159_ (.B1(_1866_),
    .Y(_1882_),
    .A1(_1864_),
    .A2(_1881_));
 sg13g2_o21ai_1 _4160_ (.B1(_1882_),
    .Y(_1883_),
    .A1(_1876_),
    .A2(_1879_));
 sg13g2_nor2b_1 _4161_ (.A(_1875_),
    .B_N(_1883_),
    .Y(_1884_));
 sg13g2_nor2_1 _4162_ (.A(_1872_),
    .B(_1884_),
    .Y(_1885_));
 sg13g2_and2_1 _4163_ (.A(_1872_),
    .B(_1884_),
    .X(_1886_));
 sg13g2_nor2_1 _4164_ (.A(_1876_),
    .B(_1882_),
    .Y(_1887_));
 sg13g2_nor2b_1 _4165_ (.A(_1887_),
    .B_N(_1879_),
    .Y(_1888_));
 sg13g2_o21ai_1 _4166_ (.B1(net1),
    .Y(_1889_),
    .A1(_1880_),
    .A2(_1888_));
 sg13g2_xor2_1 _4167_ (.B(_1883_),
    .A(_1875_),
    .X(_1890_));
 sg13g2_o21ai_1 _4168_ (.B1(_1878_),
    .Y(_1891_),
    .A1(_1856_),
    .A2(_1870_));
 sg13g2_nand2_1 _4169_ (.Y(_1892_),
    .A(_1235_),
    .B(_1891_));
 sg13g2_xnor2_1 _4170_ (.Y(_1893_),
    .A(_1890_),
    .B(_1892_));
 sg13g2_nor4_1 _4171_ (.A(_1885_),
    .B(_1886_),
    .C(_1889_),
    .D(_1893_),
    .Y(_1894_));
 sg13g2_nand2_1 _4172_ (.Y(_1895_),
    .A(_1177_),
    .B(_1234_));
 sg13g2_xor2_1 _4173_ (.B(_1786_),
    .A(_1778_),
    .X(_1896_));
 sg13g2_nand2_1 _4174_ (.Y(_1897_),
    .A(net547),
    .B(_1235_));
 sg13g2_o21ai_1 _4175_ (.B1(_1895_),
    .Y(_1898_),
    .A1(_1896_),
    .A2(_1897_));
 sg13g2_a21o_1 _4176_ (.A2(_1898_),
    .A1(_1789_),
    .B1(_1792_),
    .X(_1899_));
 sg13g2_nand3_1 _4177_ (.B(_1894_),
    .C(_1899_),
    .A(_1795_),
    .Y(_1900_));
 sg13g2_or2_1 _4178_ (.X(_1901_),
    .B(_1449_),
    .A(_1352_));
 sg13g2_nand3b_1 _4179_ (.B(_1548_),
    .C(_1620_),
    .Y(_1902_),
    .A_N(net1));
 sg13g2_nand2b_1 _4180_ (.Y(_1903_),
    .B(_1901_),
    .A_N(_1902_));
 sg13g2_a21oi_1 _4181_ (.A1(_1900_),
    .A2(_1903_),
    .Y(_0381_),
    .B1(net750));
 sg13g2_nor2_1 _4182_ (.A(_1352_),
    .B(_1720_),
    .Y(_1904_));
 sg13g2_nor2_1 _4183_ (.A(_1550_),
    .B(_1901_),
    .Y(_1905_));
 sg13g2_nor3_1 _4184_ (.A(_1352_),
    .B(_1550_),
    .C(_1720_),
    .Y(_1906_));
 sg13g2_or2_1 _4185_ (.X(_0379_),
    .B(_1906_),
    .A(_0381_));
 sg13g2_or2_1 _4186_ (.X(_0380_),
    .B(_1905_),
    .A(_0381_));
 sg13g2_nand3_1 _4187_ (.B(_1619_),
    .C(_1720_),
    .A(_1351_),
    .Y(_1907_));
 sg13g2_nand2b_1 _4188_ (.Y(_1908_),
    .B(_1907_),
    .A_N(_1902_));
 sg13g2_and2_1 _4189_ (.A(_1900_),
    .B(_1908_),
    .X(_1909_));
 sg13g2_nand2_1 _4190_ (.Y(_1910_),
    .A(_1616_),
    .B(_1905_));
 sg13g2_o21ai_1 _4191_ (.B1(_1910_),
    .Y(_0382_),
    .A1(net750),
    .A2(_1909_));
 sg13g2_o21ai_1 _4192_ (.B1(_1900_),
    .Y(_1911_),
    .A1(_1902_),
    .A2(_1904_));
 sg13g2_a21o_1 _4193_ (.A2(_1911_),
    .A1(net795),
    .B1(_1906_),
    .X(_0383_));
 sg13g2_xnor2_1 _4194_ (.Y(_1912_),
    .A(\tmds_red.n102 ),
    .B(_0891_));
 sg13g2_a21oi_1 _4195_ (.A1(net607),
    .A2(_1912_),
    .Y(_0384_),
    .B1(net750));
 sg13g2_xor2_1 _4196_ (.B(_0860_),
    .A(\tmds_red.n114 ),
    .X(_1913_));
 sg13g2_a21oi_1 _4197_ (.A1(_0891_),
    .A2(_1913_),
    .Y(_1914_),
    .B1(_0647_));
 sg13g2_o21ai_1 _4198_ (.B1(_1914_),
    .Y(_1915_),
    .A1(_0891_),
    .A2(_1913_));
 sg13g2_and2_1 _4199_ (.A(net803),
    .B(_1915_),
    .X(_0385_));
 sg13g2_xnor2_1 _4200_ (.Y(_1916_),
    .A(\tmds_red.n126 ),
    .B(_0860_));
 sg13g2_xnor2_1 _4201_ (.Y(_1917_),
    .A(_0889_),
    .B(_1916_));
 sg13g2_or2_1 _4202_ (.X(_1918_),
    .B(_0884_),
    .A(net548));
 sg13g2_inv_1 _4203_ (.Y(_1919_),
    .A(_1918_));
 sg13g2_a21oi_1 _4204_ (.A1(_0885_),
    .A2(_1916_),
    .Y(_1920_),
    .B1(_0647_));
 sg13g2_o21ai_1 _4205_ (.B1(_1920_),
    .Y(_1921_),
    .A1(_1916_),
    .A2(_1918_));
 sg13g2_a21oi_1 _4206_ (.A1(_0884_),
    .A2(_1917_),
    .Y(_1922_),
    .B1(_1921_));
 sg13g2_nor2_1 _4207_ (.A(_0648_),
    .B(_1922_),
    .Y(_0386_));
 sg13g2_nor2_1 _4208_ (.A(_0647_),
    .B(net548),
    .Y(_1923_));
 sg13g2_nor2_1 _4209_ (.A(net751),
    .B(_1923_),
    .Y(_0387_));
 sg13g2_nor2_1 _4210_ (.A(_0647_),
    .B(_0891_),
    .Y(_1924_));
 sg13g2_nor2_1 _4211_ (.A(net751),
    .B(_1924_),
    .Y(_0388_));
 sg13g2_a21oi_1 _4212_ (.A1(_0642_),
    .A2(net607),
    .Y(_0497_),
    .B1(net750));
 sg13g2_o21ai_1 _4213_ (.B1(net607),
    .Y(_1925_),
    .A1(\tmds_green.n126 ),
    .A2(_0844_));
 sg13g2_a21oi_1 _4214_ (.A1(_0844_),
    .A2(_0848_),
    .Y(_1926_),
    .B1(_1925_));
 sg13g2_nor2_1 _4215_ (.A(net750),
    .B(_1926_),
    .Y(_0498_));
 sg13g2_a21oi_1 _4216_ (.A1(\tmds_green.n100 ),
    .A2(net606),
    .Y(_0499_),
    .B1(net750));
 sg13g2_and2_1 _4217_ (.A(net607),
    .B(_0846_),
    .X(_1927_));
 sg13g2_a21oi_1 _4218_ (.A1(_0843_),
    .A2(_1927_),
    .Y(_0500_),
    .B1(net750));
 sg13g2_and2_1 _4219_ (.A(\tmds_red.dc_balancing_reg[0] ),
    .B(_0836_),
    .X(_0501_));
 sg13g2_xnor2_1 _4220_ (.Y(_1928_),
    .A(\tmds_red.n132 ),
    .B(\tmds_red.dc_balancing_reg[1] ));
 sg13g2_xnor2_1 _4221_ (.Y(_1929_),
    .A(\tmds_red.n114 ),
    .B(_1928_));
 sg13g2_inv_1 _4222_ (.Y(_1930_),
    .A(_1929_));
 sg13g2_o21ai_1 _4223_ (.B1(_0836_),
    .Y(_1931_),
    .A1(_0893_),
    .A2(_1930_));
 sg13g2_a21oi_1 _4224_ (.A1(_0893_),
    .A2(_1930_),
    .Y(_0502_),
    .B1(_1931_));
 sg13g2_xnor2_1 _4225_ (.Y(_1932_),
    .A(\tmds_red.dc_balancing_reg[2] ),
    .B(_0883_));
 sg13g2_inv_1 _4226_ (.Y(_1933_),
    .A(_1932_));
 sg13g2_nor2_1 _4227_ (.A(\tmds_red.dc_balancing_reg[1] ),
    .B(_0859_),
    .Y(_1934_));
 sg13g2_nor2b_1 _4228_ (.A(_0875_),
    .B_N(_0859_),
    .Y(_1935_));
 sg13g2_a21oi_1 _4229_ (.A1(_0859_),
    .A2(_0875_),
    .Y(_1936_),
    .B1(_1934_));
 sg13g2_nor2b_1 _4230_ (.A(_1932_),
    .B_N(_1936_),
    .Y(_1937_));
 sg13g2_xnor2_1 _4231_ (.Y(_1938_),
    .A(_1932_),
    .B(_1936_));
 sg13g2_xnor2_1 _4232_ (.Y(_1939_),
    .A(_1929_),
    .B(_1938_));
 sg13g2_nand3_1 _4233_ (.B(_1929_),
    .C(_1938_),
    .A(net548),
    .Y(_1940_));
 sg13g2_nor2_1 _4234_ (.A(_1934_),
    .B(_1935_),
    .Y(_1941_));
 sg13g2_xor2_1 _4235_ (.B(_1941_),
    .A(_1932_),
    .X(_1942_));
 sg13g2_nor2_1 _4236_ (.A(_1929_),
    .B(_1942_),
    .Y(_1943_));
 sg13g2_nor2_1 _4237_ (.A(_0855_),
    .B(_1929_),
    .Y(_1944_));
 sg13g2_nand2b_1 _4238_ (.Y(_1945_),
    .B(_1944_),
    .A_N(_1942_));
 sg13g2_inv_1 _4239_ (.Y(_1946_),
    .A(_1945_));
 sg13g2_and2_1 _4240_ (.A(_1929_),
    .B(_1942_),
    .X(_1947_));
 sg13g2_or4_1 _4241_ (.A(_0891_),
    .B(_1943_),
    .C(_1944_),
    .D(_1947_),
    .X(_1948_));
 sg13g2_o21ai_1 _4242_ (.B1(_1948_),
    .Y(_1949_),
    .A1(_0890_),
    .A2(_1945_));
 sg13g2_a21oi_1 _4243_ (.A1(_0855_),
    .A2(_1929_),
    .Y(_1950_),
    .B1(_1939_));
 sg13g2_nor2_1 _4244_ (.A(_0889_),
    .B(_1950_),
    .Y(_1951_));
 sg13g2_a221oi_1 _4245_ (.B2(_1951_),
    .C1(_1949_),
    .B1(_1940_),
    .A1(_1919_),
    .Y(_1952_),
    .A2(_1939_));
 sg13g2_nor2_1 _4246_ (.A(net570),
    .B(_1952_),
    .Y(_0503_));
 sg13g2_a21oi_1 _4247_ (.A1(_1930_),
    .A2(_1938_),
    .Y(_1953_),
    .B1(_1937_));
 sg13g2_o21ai_1 _4248_ (.B1(_0883_),
    .Y(_1954_),
    .A1(_0878_),
    .A2(_0880_));
 sg13g2_xnor2_1 _4249_ (.Y(_1955_),
    .A(_0653_),
    .B(_1954_));
 sg13g2_a21oi_1 _4250_ (.A1(_0654_),
    .A2(_0883_),
    .Y(_1956_),
    .B1(_0886_));
 sg13g2_xor2_1 _4251_ (.B(_1956_),
    .A(_1955_),
    .X(_1957_));
 sg13g2_nor2b_1 _4252_ (.A(_1953_),
    .B_N(_1957_),
    .Y(_1958_));
 sg13g2_xor2_1 _4253_ (.B(_1957_),
    .A(_1953_),
    .X(_1959_));
 sg13g2_nor2_1 _4254_ (.A(_1940_),
    .B(_1959_),
    .Y(_1960_));
 sg13g2_or2_1 _4255_ (.X(_1961_),
    .B(_1960_),
    .A(_0889_));
 sg13g2_a21oi_1 _4256_ (.A1(_1940_),
    .A2(_1959_),
    .Y(_1962_),
    .B1(_1961_));
 sg13g2_nor2_1 _4257_ (.A(_1918_),
    .B(_1959_),
    .Y(_1963_));
 sg13g2_a21o_1 _4258_ (.A2(_0883_),
    .A1(\tmds_red.dc_balancing_reg[2] ),
    .B1(_0886_),
    .X(_1964_));
 sg13g2_xnor2_1 _4259_ (.Y(_1965_),
    .A(_1955_),
    .B(_1964_));
 sg13g2_a21oi_1 _4260_ (.A1(_1933_),
    .A2(_1941_),
    .Y(_1966_),
    .B1(_1943_));
 sg13g2_and2_1 _4261_ (.A(_1965_),
    .B(_1966_),
    .X(_1967_));
 sg13g2_nor2_1 _4262_ (.A(_1965_),
    .B(_1966_),
    .Y(_1968_));
 sg13g2_nor4_1 _4263_ (.A(_0891_),
    .B(_1946_),
    .C(_1967_),
    .D(_1968_),
    .Y(_1969_));
 sg13g2_nor2_1 _4264_ (.A(_1945_),
    .B(_1965_),
    .Y(_1970_));
 sg13g2_nor2b_1 _4265_ (.A(_0890_),
    .B_N(_1970_),
    .Y(_1971_));
 sg13g2_nor4_1 _4266_ (.A(_1962_),
    .B(_1963_),
    .C(_1969_),
    .D(_1971_),
    .Y(_1972_));
 sg13g2_nor2_1 _4267_ (.A(net570),
    .B(_1972_),
    .Y(_0504_));
 sg13g2_a21oi_1 _4268_ (.A1(_1955_),
    .A2(_1956_),
    .Y(_1973_),
    .B1(_1958_));
 sg13g2_nor2b_1 _4269_ (.A(_0879_),
    .B_N(_0883_),
    .Y(_1974_));
 sg13g2_a21oi_1 _4270_ (.A1(\tmds_red.dc_balancing_reg[3] ),
    .A2(_1954_),
    .Y(_1975_),
    .B1(_1974_));
 sg13g2_xnor2_1 _4271_ (.Y(_1976_),
    .A(\tmds_red.dc_balancing_reg[4] ),
    .B(_1975_));
 sg13g2_xnor2_1 _4272_ (.Y(_1977_),
    .A(_1973_),
    .B(_1976_));
 sg13g2_nor2_1 _4273_ (.A(_1961_),
    .B(_1977_),
    .Y(_1978_));
 sg13g2_a21oi_1 _4274_ (.A1(_1955_),
    .A2(_1964_),
    .Y(_1979_),
    .B1(_1968_));
 sg13g2_a21oi_1 _4275_ (.A1(_0653_),
    .A2(_1954_),
    .Y(_1980_),
    .B1(_1974_));
 sg13g2_xnor2_1 _4276_ (.Y(_1981_),
    .A(\tmds_red.dc_balancing_reg[4] ),
    .B(_1980_));
 sg13g2_xnor2_1 _4277_ (.Y(_1982_),
    .A(_1979_),
    .B(_1981_));
 sg13g2_o21ai_1 _4278_ (.B1(_0889_),
    .Y(_1983_),
    .A1(_1970_),
    .A2(_1982_));
 sg13g2_a21oi_1 _4279_ (.A1(_1970_),
    .A2(_1982_),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_o21ai_1 _4280_ (.B1(_0884_),
    .Y(_1985_),
    .A1(_1978_),
    .A2(_1984_));
 sg13g2_nor2_1 _4281_ (.A(_1918_),
    .B(_1977_),
    .Y(_1986_));
 sg13g2_a21oi_1 _4282_ (.A1(_0885_),
    .A2(_1982_),
    .Y(_1987_),
    .B1(_1986_));
 sg13g2_a21oi_1 _4283_ (.A1(_1985_),
    .A2(_1987_),
    .Y(_0505_),
    .B1(net570));
 sg13g2_or4_1 _4284_ (.A(\tmds_blue.dc_balancing_reg[0] ),
    .B(\tmds_blue.dc_balancing_reg[1] ),
    .C(\tmds_blue.dc_balancing_reg[3] ),
    .D(\tmds_blue.dc_balancing_reg[2] ),
    .X(_1988_));
 sg13g2_nand2b_2 _4285_ (.Y(_1989_),
    .B(_0644_),
    .A_N(_1988_));
 sg13g2_nand3_1 _4286_ (.B(_0644_),
    .C(_1988_),
    .A(\tmds_blue.n193 ),
    .Y(_1990_));
 sg13g2_o21ai_1 _4287_ (.B1(_1990_),
    .Y(_1991_),
    .A1(\tmds_blue.n193 ),
    .A2(_0644_));
 sg13g2_xnor2_1 _4288_ (.Y(_1992_),
    .A(_0643_),
    .B(_1991_));
 sg13g2_nand2_1 _4289_ (.Y(_1993_),
    .A(_1989_),
    .B(_1992_));
 sg13g2_o21ai_1 _4290_ (.B1(net797),
    .Y(_1994_),
    .A1(net607),
    .A2(hsync));
 sg13g2_a21oi_1 _4291_ (.A1(net606),
    .A2(_1993_),
    .Y(_0610_),
    .B1(_1994_));
 sg13g2_nand2_1 _4292_ (.Y(_1995_),
    .A(_0643_),
    .B(\tmds_blue.n193 ));
 sg13g2_xnor2_1 _4293_ (.Y(_1996_),
    .A(net604),
    .B(\tmds_blue.n193 ));
 sg13g2_o21ai_1 _4294_ (.B1(net606),
    .Y(_1997_),
    .A1(_1988_),
    .A2(_1996_));
 sg13g2_nor2_2 _4295_ (.A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_1997_),
    .Y(_1998_));
 sg13g2_nor2_1 _4296_ (.A(_1994_),
    .B(_1998_),
    .Y(_0611_));
 sg13g2_nor2b_1 _4297_ (.A(net606),
    .B_N(hsync),
    .Y(_1999_));
 sg13g2_nand2b_1 _4298_ (.Y(_2000_),
    .B(net797),
    .A_N(_1999_));
 sg13g2_nor2_1 _4299_ (.A(_1998_),
    .B(_2000_),
    .Y(_0612_));
 sg13g2_xnor2_1 _4300_ (.Y(_2001_),
    .A(\tmds_blue.n126 ),
    .B(_1996_));
 sg13g2_nor2b_2 _4301_ (.A(_1991_),
    .B_N(_1989_),
    .Y(_2002_));
 sg13g2_inv_1 _4302_ (.Y(_2003_),
    .A(_2002_));
 sg13g2_nor2_2 _4303_ (.A(net604),
    .B(_1989_),
    .Y(_2004_));
 sg13g2_o21ai_1 _4304_ (.B1(net606),
    .Y(_2005_),
    .A1(_2002_),
    .A2(_2004_));
 sg13g2_or3_1 _4305_ (.A(_0647_),
    .B(_2002_),
    .C(_2004_),
    .X(_2006_));
 sg13g2_mux2_1 _4306_ (.A0(_2005_),
    .A1(_2006_),
    .S(_2001_),
    .X(_2007_));
 sg13g2_nor2b_1 _4307_ (.A(_2000_),
    .B_N(_2007_),
    .Y(_0615_));
 sg13g2_xor2_1 _4308_ (.B(\tmds_blue.n132 ),
    .A(net605),
    .X(_2008_));
 sg13g2_xnor2_1 _4309_ (.Y(_2009_),
    .A(_2001_),
    .B(_2008_));
 sg13g2_nand2b_1 _4310_ (.Y(_2010_),
    .B(_2009_),
    .A_N(_2006_));
 sg13g2_nor2_1 _4311_ (.A(_2005_),
    .B(_2009_),
    .Y(_2011_));
 sg13g2_nor2_1 _4312_ (.A(_1999_),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_1 _4313_ (.A1(_2010_),
    .A2(_2012_),
    .Y(_0616_),
    .B1(net749));
 sg13g2_a21oi_1 _4314_ (.A1(net605),
    .A2(net607),
    .Y(_0617_),
    .B1(_2000_));
 sg13g2_o21ai_1 _4315_ (.B1(\tmds_blue.vsync ),
    .Y(_2013_),
    .A1(net606),
    .A2(hsync));
 sg13g2_o21ai_1 _4316_ (.B1(_2013_),
    .Y(_2014_),
    .A1(\tmds_blue.vsync ),
    .A2(_1999_));
 sg13g2_and3_1 _4317_ (.X(_0618_),
    .A(net797),
    .B(_2005_),
    .C(_2014_));
 sg13g2_nand2b_1 _4318_ (.Y(_2015_),
    .B(\tmds_green.dc_balancing_reg[1] ),
    .A_N(net601));
 sg13g2_nand2b_2 _4319_ (.Y(_2016_),
    .B(net601),
    .A_N(\tmds_green.dc_balancing_reg[1] ));
 sg13g2_nand3_1 _4320_ (.B(_2015_),
    .C(_2016_),
    .A(net602),
    .Y(_2017_));
 sg13g2_a21o_1 _4321_ (.A2(_2016_),
    .A1(_2015_),
    .B1(net602),
    .X(_2018_));
 sg13g2_and2_1 _4322_ (.A(_2017_),
    .B(_2018_),
    .X(_2019_));
 sg13g2_xnor2_1 _4323_ (.Y(_2020_),
    .A(_0642_),
    .B(_2019_));
 sg13g2_nor2_1 _4324_ (.A(net569),
    .B(_2020_),
    .Y(_0619_));
 sg13g2_nor2_1 _4325_ (.A(net601),
    .B(\tmds_green.n126 ),
    .Y(_2021_));
 sg13g2_nor3_1 _4326_ (.A(net603),
    .B(net601),
    .C(\tmds_green.n126 ),
    .Y(_2022_));
 sg13g2_nand2_1 _4327_ (.Y(_2023_),
    .A(net601),
    .B(\tmds_green.n126 ));
 sg13g2_nand3_1 _4328_ (.B(\tmds_green.n132 ),
    .C(\tmds_green.n126 ),
    .A(net603),
    .Y(_2024_));
 sg13g2_nor2_1 _4329_ (.A(net602),
    .B(_2021_),
    .Y(_2025_));
 sg13g2_nand2_1 _4330_ (.Y(_2026_),
    .A(net602),
    .B(_2023_));
 sg13g2_nand2b_2 _4331_ (.Y(_2027_),
    .B(_2024_),
    .A_N(_2022_));
 sg13g2_nand2b_1 _4332_ (.Y(_2028_),
    .B(_2027_),
    .A_N(\tmds_green.dc_balancing_reg[2] ));
 sg13g2_xor2_1 _4333_ (.B(_2027_),
    .A(\tmds_green.dc_balancing_reg[2] ),
    .X(_2029_));
 sg13g2_and2_1 _4334_ (.A(_2016_),
    .B(_2029_),
    .X(_2030_));
 sg13g2_nand2_1 _4335_ (.Y(_2031_),
    .A(_2016_),
    .B(_2029_));
 sg13g2_xor2_1 _4336_ (.B(_2029_),
    .A(_2016_),
    .X(_2032_));
 sg13g2_o21ai_1 _4337_ (.B1(_0841_),
    .Y(_2033_),
    .A1(\tmds_green.dc_balancing_reg[1] ),
    .A2(_0842_));
 sg13g2_nor2b_1 _4338_ (.A(_2033_),
    .B_N(_2029_),
    .Y(_2034_));
 sg13g2_nand2b_1 _4339_ (.Y(_2035_),
    .B(_2033_),
    .A_N(_2029_));
 sg13g2_nor2b_1 _4340_ (.A(_2034_),
    .B_N(_2035_),
    .Y(_2036_));
 sg13g2_xnor2_1 _4341_ (.Y(_2037_),
    .A(_2017_),
    .B(_2036_));
 sg13g2_nand2_1 _4342_ (.Y(_2038_),
    .A(_0847_),
    .B(_2037_));
 sg13g2_o21ai_1 _4343_ (.B1(_2038_),
    .Y(_2039_),
    .A1(_0847_),
    .A2(_2032_));
 sg13g2_xnor2_1 _4344_ (.Y(_2040_),
    .A(_0844_),
    .B(_2039_));
 sg13g2_nor2_1 _4345_ (.A(net569),
    .B(_2040_),
    .Y(_0620_));
 sg13g2_nor2_1 _4346_ (.A(_2018_),
    .B(_2029_),
    .Y(_2041_));
 sg13g2_xnor2_1 _4347_ (.Y(_2042_),
    .A(_0641_),
    .B(_2027_));
 sg13g2_inv_1 _4348_ (.Y(_2043_),
    .A(_2042_));
 sg13g2_nand2_1 _4349_ (.Y(_2044_),
    .A(_2026_),
    .B(_2028_));
 sg13g2_nor2_1 _4350_ (.A(_2042_),
    .B(_2044_),
    .Y(_2045_));
 sg13g2_xnor2_1 _4351_ (.Y(_2046_),
    .A(_2043_),
    .B(_2044_));
 sg13g2_a21oi_1 _4352_ (.A1(_2019_),
    .A2(_2035_),
    .Y(_2047_),
    .B1(_2034_));
 sg13g2_inv_1 _4353_ (.Y(_2048_),
    .A(_2047_));
 sg13g2_xor2_1 _4354_ (.B(_2047_),
    .A(_2046_),
    .X(_2049_));
 sg13g2_nor3_1 _4355_ (.A(_2018_),
    .B(_2029_),
    .C(_2049_),
    .Y(_2050_));
 sg13g2_a21oi_1 _4356_ (.A1(_2046_),
    .A2(_2048_),
    .Y(_2051_),
    .B1(_2045_));
 sg13g2_a21oi_1 _4357_ (.A1(\tmds_green.dc_balancing_reg[3] ),
    .A2(_2024_),
    .Y(_2052_),
    .B1(_2022_));
 sg13g2_xnor2_1 _4358_ (.Y(_2053_),
    .A(\tmds_green.dc_balancing_reg[4] ),
    .B(_2052_));
 sg13g2_xnor2_1 _4359_ (.Y(_2054_),
    .A(_2051_),
    .B(_2053_));
 sg13g2_xnor2_1 _4360_ (.Y(_2055_),
    .A(_2041_),
    .B(_2049_));
 sg13g2_nor2b_1 _4361_ (.A(_2025_),
    .B_N(_2028_),
    .Y(_2056_));
 sg13g2_nor2_1 _4362_ (.A(_2043_),
    .B(_2056_),
    .Y(_2057_));
 sg13g2_xnor2_1 _4363_ (.Y(_2058_),
    .A(_2042_),
    .B(_2056_));
 sg13g2_xnor2_1 _4364_ (.Y(_2059_),
    .A(_2031_),
    .B(_2058_));
 sg13g2_nand2b_1 _4365_ (.Y(_2060_),
    .B(_2059_),
    .A_N(_0847_));
 sg13g2_a21oi_1 _4366_ (.A1(_0847_),
    .A2(_2055_),
    .Y(_2061_),
    .B1(_0840_));
 sg13g2_a21oi_1 _4367_ (.A1(_2060_),
    .A2(_2061_),
    .Y(_0621_),
    .B1(net570));
 sg13g2_xnor2_1 _4368_ (.Y(_2062_),
    .A(_2050_),
    .B(_2054_));
 sg13g2_nand2_1 _4369_ (.Y(_2063_),
    .A(_0847_),
    .B(_2062_));
 sg13g2_nand2b_1 _4370_ (.Y(_2064_),
    .B(_2015_),
    .A_N(_2029_));
 sg13g2_nand4_1 _4371_ (.B(_2031_),
    .C(_2058_),
    .A(net602),
    .Y(_2065_),
    .D(_2064_));
 sg13g2_a221oi_1 _4372_ (.B2(net603),
    .C1(_2030_),
    .B1(_2064_),
    .A1(_2043_),
    .Y(_2066_),
    .A2(_2056_));
 sg13g2_nor2_1 _4373_ (.A(_2057_),
    .B(_2066_),
    .Y(_2067_));
 sg13g2_o21ai_1 _4374_ (.B1(_2024_),
    .Y(_2068_),
    .A1(_0641_),
    .A2(_2022_));
 sg13g2_xnor2_1 _4375_ (.Y(_2069_),
    .A(\tmds_green.dc_balancing_reg[4] ),
    .B(_2068_));
 sg13g2_xnor2_1 _4376_ (.Y(_2070_),
    .A(_2067_),
    .B(_2069_));
 sg13g2_a21oi_1 _4377_ (.A1(_2065_),
    .A2(_2070_),
    .Y(_2071_),
    .B1(_0847_));
 sg13g2_nor2_1 _4378_ (.A(_0840_),
    .B(_2071_),
    .Y(_2072_));
 sg13g2_a21oi_1 _4379_ (.A1(_2063_),
    .A2(_2072_),
    .Y(_0622_),
    .B1(net570));
 sg13g2_nor3_1 _4380_ (.A(net749),
    .B(\clockdiv.q0 ),
    .C(net406),
    .Y(_0623_));
 sg13g2_xor2_1 _4381_ (.B(\tmds_blue.dc_balancing_reg[1] ),
    .A(\tmds_blue.n193 ),
    .X(_2073_));
 sg13g2_xnor2_1 _4382_ (.Y(_2074_),
    .A(\tmds_blue.n132 ),
    .B(_2073_));
 sg13g2_o21ai_1 _4383_ (.B1(_0836_),
    .Y(_2075_),
    .A1(_1993_),
    .A2(_2074_));
 sg13g2_a21oi_1 _4384_ (.A1(_1993_),
    .A2(_2074_),
    .Y(_0624_),
    .B1(_2075_));
 sg13g2_xor2_1 _4385_ (.B(\tmds_blue.n193 ),
    .A(\tmds_blue.n132 ),
    .X(_2076_));
 sg13g2_and2_1 _4386_ (.A(\tmds_blue.n126 ),
    .B(\tmds_blue.n132 ),
    .X(_2077_));
 sg13g2_nor3_1 _4387_ (.A(net604),
    .B(_2001_),
    .C(_2077_),
    .Y(_2078_));
 sg13g2_a21oi_1 _4388_ (.A1(_1995_),
    .A2(_2077_),
    .Y(_2079_),
    .B1(_2078_));
 sg13g2_nor2_2 _4389_ (.A(_2076_),
    .B(_2079_),
    .Y(_2080_));
 sg13g2_nand2b_1 _4390_ (.Y(_2081_),
    .B(_2080_),
    .A_N(\tmds_blue.dc_balancing_reg[2] ));
 sg13g2_xnor2_1 _4391_ (.Y(_2082_),
    .A(\tmds_blue.dc_balancing_reg[2] ),
    .B(_2080_));
 sg13g2_nand2b_1 _4392_ (.Y(_2083_),
    .B(_2076_),
    .A_N(_2079_));
 sg13g2_o21ai_1 _4393_ (.B1(_2083_),
    .Y(_2084_),
    .A1(\tmds_blue.dc_balancing_reg[1] ),
    .A2(_2076_));
 sg13g2_nor2_1 _4394_ (.A(_2082_),
    .B(_2084_),
    .Y(_2085_));
 sg13g2_xor2_1 _4395_ (.B(_2084_),
    .A(_2082_),
    .X(_2086_));
 sg13g2_and2_1 _4396_ (.A(_2074_),
    .B(_2086_),
    .X(_2087_));
 sg13g2_xnor2_1 _4397_ (.Y(_2088_),
    .A(_2074_),
    .B(_2086_));
 sg13g2_o21ai_1 _4398_ (.B1(_2083_),
    .Y(_2089_),
    .A1(_0645_),
    .A2(_2076_));
 sg13g2_inv_1 _4399_ (.Y(_2090_),
    .A(_2089_));
 sg13g2_xor2_1 _4400_ (.B(_2089_),
    .A(_2082_),
    .X(_2091_));
 sg13g2_nand2b_1 _4401_ (.Y(_2092_),
    .B(_2074_),
    .A_N(_2091_));
 sg13g2_nor2_1 _4402_ (.A(net604),
    .B(_2074_),
    .Y(_2093_));
 sg13g2_xnor2_1 _4403_ (.Y(_2094_),
    .A(_2074_),
    .B(_2091_));
 sg13g2_nor3_1 _4404_ (.A(_2004_),
    .B(_2093_),
    .C(_2094_),
    .Y(_2095_));
 sg13g2_nor2b_1 _4405_ (.A(_2091_),
    .B_N(_2093_),
    .Y(_2096_));
 sg13g2_inv_1 _4406_ (.Y(_2097_),
    .A(_2096_));
 sg13g2_a221oi_1 _4407_ (.B2(_1989_),
    .C1(_2095_),
    .B1(_2096_),
    .A1(_2004_),
    .Y(_2098_),
    .A2(_2088_));
 sg13g2_nor2_1 _4408_ (.A(_2002_),
    .B(_2098_),
    .Y(_2099_));
 sg13g2_a21oi_1 _4409_ (.A1(net604),
    .A2(_2074_),
    .Y(_2100_),
    .B1(_2088_));
 sg13g2_and2_1 _4410_ (.A(net605),
    .B(_2087_),
    .X(_2101_));
 sg13g2_inv_1 _4411_ (.Y(_2102_),
    .A(_2101_));
 sg13g2_nor3_1 _4412_ (.A(_2003_),
    .B(_2100_),
    .C(_2101_),
    .Y(_2103_));
 sg13g2_nor3_1 _4413_ (.A(net571),
    .B(_2099_),
    .C(_2103_),
    .Y(_0625_));
 sg13g2_nor2_1 _4414_ (.A(_2085_),
    .B(_2087_),
    .Y(_2104_));
 sg13g2_nand2_1 _4415_ (.Y(_2105_),
    .A(net604),
    .B(_2077_));
 sg13g2_nand2_1 _4416_ (.Y(_2106_),
    .A(\tmds_blue.n193 ),
    .B(_2105_));
 sg13g2_inv_1 _4417_ (.Y(_2107_),
    .A(_2106_));
 sg13g2_o21ai_1 _4418_ (.B1(_2081_),
    .Y(_2108_),
    .A1(_2080_),
    .A2(_2107_));
 sg13g2_xnor2_1 _4419_ (.Y(_2109_),
    .A(\tmds_blue.dc_balancing_reg[3] ),
    .B(_2080_));
 sg13g2_nand2b_1 _4420_ (.Y(_2110_),
    .B(_2109_),
    .A_N(_2108_));
 sg13g2_xnor2_1 _4421_ (.Y(_2111_),
    .A(_2108_),
    .B(_2109_));
 sg13g2_o21ai_1 _4422_ (.B1(_2111_),
    .Y(_2112_),
    .A1(_2085_),
    .A2(_2087_));
 sg13g2_xnor2_1 _4423_ (.Y(_2113_),
    .A(_2104_),
    .B(_2111_));
 sg13g2_o21ai_1 _4424_ (.B1(_2092_),
    .Y(_2114_),
    .A1(_2082_),
    .A2(_2090_));
 sg13g2_inv_1 _4425_ (.Y(_2115_),
    .A(_2114_));
 sg13g2_nand3_1 _4426_ (.B(_2106_),
    .C(_2109_),
    .A(_2081_),
    .Y(_2116_));
 sg13g2_a21o_1 _4427_ (.A2(_2106_),
    .A1(_2081_),
    .B1(_2109_),
    .X(_2117_));
 sg13g2_nand2_1 _4428_ (.Y(_2118_),
    .A(_2116_),
    .B(_2117_));
 sg13g2_xor2_1 _4429_ (.B(_2118_),
    .A(_2114_),
    .X(_2119_));
 sg13g2_nor3_1 _4430_ (.A(_0643_),
    .B(_1989_),
    .C(_2119_),
    .Y(_2120_));
 sg13g2_a21oi_1 _4431_ (.A1(_2004_),
    .A2(_2113_),
    .Y(_2121_),
    .B1(_2120_));
 sg13g2_xnor2_1 _4432_ (.Y(_2122_),
    .A(_2097_),
    .B(_2119_));
 sg13g2_nand2_1 _4433_ (.Y(_2123_),
    .A(_2101_),
    .B(_2111_));
 sg13g2_a21oi_1 _4434_ (.A1(_2102_),
    .A2(_2113_),
    .Y(_2124_),
    .B1(_1991_));
 sg13g2_a22oi_1 _4435_ (.Y(_2125_),
    .B1(_2123_),
    .B2(_2124_),
    .A2(_2122_),
    .A1(_1991_));
 sg13g2_nand2_1 _4436_ (.Y(_2126_),
    .A(_1989_),
    .B(_2125_));
 sg13g2_a21oi_1 _4437_ (.A1(_2121_),
    .A2(_2126_),
    .Y(_0626_),
    .B1(net571));
 sg13g2_o21ai_1 _4438_ (.B1(_2116_),
    .Y(_2127_),
    .A1(_2115_),
    .A2(_2118_));
 sg13g2_nand3_1 _4439_ (.B(\tmds_blue.n193 ),
    .C(_2077_),
    .A(net604),
    .Y(_2128_));
 sg13g2_o21ai_1 _4440_ (.B1(_2128_),
    .Y(_2129_),
    .A1(\tmds_blue.dc_balancing_reg[3] ),
    .A2(_2080_));
 sg13g2_xnor2_1 _4441_ (.Y(_2130_),
    .A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_2129_));
 sg13g2_xnor2_1 _4442_ (.Y(_2131_),
    .A(_2127_),
    .B(_2130_));
 sg13g2_o21ai_1 _4443_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2097_),
    .A2(_2119_));
 sg13g2_o21ai_1 _4444_ (.B1(_2128_),
    .Y(_2133_),
    .A1(_0646_),
    .A2(_2080_));
 sg13g2_xnor2_1 _4445_ (.Y(_2134_),
    .A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_2133_));
 sg13g2_a21oi_1 _4446_ (.A1(_2110_),
    .A2(_2112_),
    .Y(_2135_),
    .B1(_2134_));
 sg13g2_nand3_1 _4447_ (.B(_2112_),
    .C(_2134_),
    .A(_2110_),
    .Y(_2136_));
 sg13g2_nand3b_1 _4448_ (.B(_2123_),
    .C(_2136_),
    .Y(_2137_),
    .A_N(_1991_));
 sg13g2_o21ai_1 _4449_ (.B1(_1989_),
    .Y(_2138_),
    .A1(_2135_),
    .A2(_2137_));
 sg13g2_a21o_1 _4450_ (.A2(_2132_),
    .A1(_1991_),
    .B1(_2138_),
    .X(_2139_));
 sg13g2_a21oi_1 _4451_ (.A1(_2121_),
    .A2(_2139_),
    .Y(_0627_),
    .B1(net571));
 sg13g2_nor2_1 _4452_ (.A(net680),
    .B(net731),
    .Y(_0007_));
 sg13g2_nor2_1 _4453_ (.A(net682),
    .B(net733),
    .Y(_0008_));
 sg13g2_nor2_1 _4454_ (.A(net679),
    .B(net730),
    .Y(_0009_));
 sg13g2_nor2_1 _4455_ (.A(_0642_),
    .B(net569),
    .Y(_0272_));
 sg13g2_nor2_1 _4456_ (.A(net569),
    .B(_0894_),
    .Y(_0277_));
 sg13g2_nor2_1 _4457_ (.A(net657),
    .B(net708),
    .Y(_0010_));
 sg13g2_nor2_1 _4458_ (.A(net651),
    .B(net707),
    .Y(_0011_));
 sg13g2_nor2_1 _4459_ (.A(net656),
    .B(net702),
    .Y(_0012_));
 sg13g2_nor2_1 _4460_ (.A(net651),
    .B(net702),
    .Y(_0013_));
 sg13g2_nor2_1 _4461_ (.A(net663),
    .B(net714),
    .Y(_0014_));
 sg13g2_nor2_1 _4462_ (.A(net659),
    .B(net710),
    .Y(_0015_));
 sg13g2_nor2_1 _4463_ (.A(net668),
    .B(net720),
    .Y(_0016_));
 sg13g2_nor2_1 _4464_ (.A(net655),
    .B(net706),
    .Y(_0017_));
 sg13g2_nor2_1 _4465_ (.A(net675),
    .B(net725),
    .Y(_0018_));
 sg13g2_nor2_1 _4466_ (.A(net674),
    .B(net725),
    .Y(_0019_));
 sg13g2_nor2_1 _4467_ (.A(net675),
    .B(net727),
    .Y(_0020_));
 sg13g2_nor2_1 _4468_ (.A(net674),
    .B(net726),
    .Y(_0021_));
 sg13g2_nor2_1 _4469_ (.A(net661),
    .B(net712),
    .Y(_0022_));
 sg13g2_nor2_1 _4470_ (.A(net664),
    .B(net715),
    .Y(_0023_));
 sg13g2_nor2_1 _4471_ (.A(net662),
    .B(net713),
    .Y(_0024_));
 sg13g2_nor2_1 _4472_ (.A(net664),
    .B(net715),
    .Y(_0025_));
 sg13g2_nor2_1 _4473_ (.A(net661),
    .B(net712),
    .Y(_0026_));
 sg13g2_nor2_1 _4474_ (.A(net659),
    .B(net710),
    .Y(_0027_));
 sg13g2_nor2_1 _4475_ (.A(net668),
    .B(net720),
    .Y(_0028_));
 sg13g2_nor2_1 _4476_ (.A(net653),
    .B(net704),
    .Y(_0029_));
 sg13g2_nor2_1 _4477_ (.A(net661),
    .B(net712),
    .Y(_0030_));
 sg13g2_nor2_1 _4478_ (.A(net665),
    .B(net716),
    .Y(_0031_));
 sg13g2_nor2_1 _4479_ (.A(net662),
    .B(net713),
    .Y(_0032_));
 sg13g2_nor2_1 _4480_ (.A(net664),
    .B(net715),
    .Y(_0033_));
 sg13g2_nor2_1 _4481_ (.A(net670),
    .B(net721),
    .Y(_0034_));
 sg13g2_nor2_1 _4482_ (.A(net670),
    .B(net721),
    .Y(_0035_));
 sg13g2_nor2_1 _4483_ (.A(net670),
    .B(net721),
    .Y(_0036_));
 sg13g2_nor2_1 _4484_ (.A(net670),
    .B(net721),
    .Y(_0037_));
 sg13g2_nor2_1 _4485_ (.A(net686),
    .B(net737),
    .Y(_0038_));
 sg13g2_nor2_1 _4486_ (.A(net685),
    .B(net736),
    .Y(_0039_));
 sg13g2_nor2_1 _4487_ (.A(net685),
    .B(net736),
    .Y(_0040_));
 sg13g2_nor2_1 _4488_ (.A(net684),
    .B(net735),
    .Y(_0041_));
 sg13g2_nor2_1 _4489_ (.A(net653),
    .B(net704),
    .Y(_0042_));
 sg13g2_nor2_1 _4490_ (.A(net652),
    .B(net703),
    .Y(_0043_));
 sg13g2_nor2_1 _4491_ (.A(net653),
    .B(net704),
    .Y(_0044_));
 sg13g2_nor2_1 _4492_ (.A(net652),
    .B(net703),
    .Y(_0045_));
 sg13g2_nor2_1 _4493_ (.A(net651),
    .B(net702),
    .Y(_0046_));
 sg13g2_nor2_1 _4494_ (.A(net651),
    .B(net702),
    .Y(_0047_));
 sg13g2_nor2_1 _4495_ (.A(net652),
    .B(net703),
    .Y(_0048_));
 sg13g2_nor2_1 _4496_ (.A(net651),
    .B(net702),
    .Y(_0049_));
 sg13g2_nor2_1 _4497_ (.A(net651),
    .B(net702),
    .Y(_0050_));
 sg13g2_nor2_1 _4498_ (.A(net652),
    .B(net703),
    .Y(_0051_));
 sg13g2_nor2_1 _4499_ (.A(net652),
    .B(net703),
    .Y(_0052_));
 sg13g2_nor2_1 _4500_ (.A(net652),
    .B(net703),
    .Y(_0053_));
 sg13g2_nor2_1 _4501_ (.A(net651),
    .B(net702),
    .Y(_0054_));
 sg13g2_nor2_1 _4502_ (.A(net656),
    .B(net707),
    .Y(_0055_));
 sg13g2_nor2_1 _4503_ (.A(net652),
    .B(net703),
    .Y(_0056_));
 sg13g2_nor2_1 _4504_ (.A(net651),
    .B(net702),
    .Y(_0057_));
 sg13g2_nor2_1 _4505_ (.A(net663),
    .B(net724),
    .Y(_0058_));
 sg13g2_nor2_1 _4506_ (.A(net659),
    .B(net710),
    .Y(_0059_));
 sg13g2_nor2_1 _4507_ (.A(net668),
    .B(net720),
    .Y(_0060_));
 sg13g2_nor2_1 _4508_ (.A(net655),
    .B(net706),
    .Y(_0061_));
 sg13g2_nor2_1 _4509_ (.A(net675),
    .B(net725),
    .Y(_0062_));
 sg13g2_nor2_1 _4510_ (.A(net674),
    .B(net726),
    .Y(_0063_));
 sg13g2_nor2_1 _4511_ (.A(net675),
    .B(net725),
    .Y(_0064_));
 sg13g2_nor2_1 _4512_ (.A(net674),
    .B(net726),
    .Y(_0065_));
 sg13g2_nor2_1 _4513_ (.A(net675),
    .B(net725),
    .Y(_0066_));
 sg13g2_nor2_1 _4514_ (.A(net674),
    .B(net727),
    .Y(_0067_));
 sg13g2_nor2_1 _4515_ (.A(net675),
    .B(net725),
    .Y(_0068_));
 sg13g2_nor2_1 _4516_ (.A(net674),
    .B(net725),
    .Y(_0069_));
 sg13g2_nor2_1 _4517_ (.A(net675),
    .B(net725),
    .Y(_0070_));
 sg13g2_nor2_1 _4518_ (.A(net674),
    .B(net726),
    .Y(_0071_));
 sg13g2_nor2_1 _4519_ (.A(net676),
    .B(net728),
    .Y(_0072_));
 sg13g2_nor2_1 _4520_ (.A(net678),
    .B(net726),
    .Y(_0073_));
 sg13g2_nor2_1 _4521_ (.A(net658),
    .B(net709),
    .Y(_0074_));
 sg13g2_nor2_1 _4522_ (.A(net657),
    .B(net708),
    .Y(_0075_));
 sg13g2_nor2_1 _4523_ (.A(net675),
    .B(net709),
    .Y(_0076_));
 sg13g2_nor2_1 _4524_ (.A(net658),
    .B(net708),
    .Y(_0077_));
 sg13g2_nor2_1 _4525_ (.A(net658),
    .B(net709),
    .Y(_0078_));
 sg13g2_nor2_1 _4526_ (.A(net657),
    .B(net708),
    .Y(_0079_));
 sg13g2_nor2_1 _4527_ (.A(net658),
    .B(net709),
    .Y(_0080_));
 sg13g2_nor2_1 _4528_ (.A(net657),
    .B(net708),
    .Y(_0081_));
 sg13g2_nor2_1 _4529_ (.A(net658),
    .B(net709),
    .Y(_0082_));
 sg13g2_nor2_1 _4530_ (.A(net657),
    .B(net708),
    .Y(_0083_));
 sg13g2_nor2_1 _4531_ (.A(net657),
    .B(net708),
    .Y(_0084_));
 sg13g2_nor2_1 _4532_ (.A(net657),
    .B(net708),
    .Y(_0085_));
 sg13g2_nor2_1 _4533_ (.A(net660),
    .B(net711),
    .Y(_0086_));
 sg13g2_nor2_1 _4534_ (.A(net660),
    .B(net711),
    .Y(_0087_));
 sg13g2_nor2_1 _4535_ (.A(net659),
    .B(net710),
    .Y(_0088_));
 sg13g2_nor2_1 _4536_ (.A(net657),
    .B(net709),
    .Y(_0089_));
 sg13g2_nor2_1 _4537_ (.A(net679),
    .B(net726),
    .Y(_0090_));
 sg13g2_nor2_1 _4538_ (.A(net679),
    .B(net730),
    .Y(_0091_));
 sg13g2_nor2_1 _4539_ (.A(net680),
    .B(net726),
    .Y(_0092_));
 sg13g2_nor2_1 _4540_ (.A(net679),
    .B(net730),
    .Y(_0093_));
 sg13g2_nor2_1 _4541_ (.A(net674),
    .B(net726),
    .Y(_0094_));
 sg13g2_nor2_1 _4542_ (.A(net679),
    .B(net730),
    .Y(_0095_));
 sg13g2_nor2_1 _4543_ (.A(net680),
    .B(net731),
    .Y(_0096_));
 sg13g2_nor2_1 _4544_ (.A(net679),
    .B(net730),
    .Y(_0097_));
 sg13g2_nor2_1 _4545_ (.A(net661),
    .B(net712),
    .Y(_0098_));
 sg13g2_nor2_1 _4546_ (.A(net655),
    .B(net706),
    .Y(_0099_));
 sg13g2_nor2_1 _4547_ (.A(net668),
    .B(net720),
    .Y(_0100_));
 sg13g2_nor2_1 _4548_ (.A(net655),
    .B(net706),
    .Y(_0101_));
 sg13g2_nor2_1 _4549_ (.A(net679),
    .B(net730),
    .Y(_0102_));
 sg13g2_nor2_1 _4550_ (.A(net680),
    .B(net731),
    .Y(_0103_));
 sg13g2_nor2_1 _4551_ (.A(net680),
    .B(net730),
    .Y(_0104_));
 sg13g2_nor2_1 _4552_ (.A(net680),
    .B(net731),
    .Y(_0105_));
 sg13g2_nor2_1 _4553_ (.A(net682),
    .B(net733),
    .Y(_0106_));
 sg13g2_nor2_1 _4554_ (.A(net682),
    .B(net733),
    .Y(_0107_));
 sg13g2_nor2_1 _4555_ (.A(net682),
    .B(net733),
    .Y(_0108_));
 sg13g2_nor2_1 _4556_ (.A(net682),
    .B(net733),
    .Y(_0109_));
 sg13g2_nor2_1 _4557_ (.A(net681),
    .B(net732),
    .Y(_0110_));
 sg13g2_nor2_1 _4558_ (.A(net689),
    .B(net741),
    .Y(_0111_));
 sg13g2_nor2_1 _4559_ (.A(net682),
    .B(net733),
    .Y(_0112_));
 sg13g2_nor2_1 _4560_ (.A(net681),
    .B(net732),
    .Y(_0113_));
 sg13g2_nor2_1 _4561_ (.A(net681),
    .B(net732),
    .Y(_0114_));
 sg13g2_nor2_1 _4562_ (.A(net681),
    .B(net732),
    .Y(_0115_));
 sg13g2_nor2_1 _4563_ (.A(net682),
    .B(net733),
    .Y(_0116_));
 sg13g2_nor2_1 _4564_ (.A(net681),
    .B(net732),
    .Y(_0117_));
 sg13g2_nor2_1 _4565_ (.A(net681),
    .B(net732),
    .Y(_0118_));
 sg13g2_nor2_1 _4566_ (.A(net683),
    .B(net732),
    .Y(_0119_));
 sg13g2_nor2_1 _4567_ (.A(net681),
    .B(net732),
    .Y(_0120_));
 sg13g2_nor2_1 _4568_ (.A(net681),
    .B(net734),
    .Y(_0121_));
 sg13g2_nor2_1 _4569_ (.A(net676),
    .B(net728),
    .Y(_0122_));
 sg13g2_nor2_1 _4570_ (.A(net684),
    .B(net735),
    .Y(_0123_));
 sg13g2_nor2_1 _4571_ (.A(net677),
    .B(net729),
    .Y(_0124_));
 sg13g2_nor2_1 _4572_ (.A(net685),
    .B(net736),
    .Y(_0125_));
 sg13g2_nor2_1 _4573_ (.A(net676),
    .B(net728),
    .Y(_0126_));
 sg13g2_nor2_1 _4574_ (.A(net685),
    .B(net736),
    .Y(_0127_));
 sg13g2_nor2_1 _4575_ (.A(net676),
    .B(net728),
    .Y(_0128_));
 sg13g2_nor2_1 _4576_ (.A(net685),
    .B(net736),
    .Y(_0129_));
 sg13g2_nor2_1 _4577_ (.A(net661),
    .B(net712),
    .Y(_0130_));
 sg13g2_nor2_1 _4578_ (.A(net664),
    .B(net715),
    .Y(_0131_));
 sg13g2_nor2_1 _4579_ (.A(net663),
    .B(net714),
    .Y(_0132_));
 sg13g2_nor2_1 _4580_ (.A(net666),
    .B(net717),
    .Y(_0133_));
 sg13g2_nor2_1 _4581_ (.A(net676),
    .B(net728),
    .Y(_0134_));
 sg13g2_nor2_1 _4582_ (.A(net677),
    .B(net728),
    .Y(_0135_));
 sg13g2_nor2_1 _4583_ (.A(net677),
    .B(net729),
    .Y(_0136_));
 sg13g2_nor2_1 _4584_ (.A(net677),
    .B(net729),
    .Y(_0137_));
 sg13g2_nor2_1 _4585_ (.A(net676),
    .B(net728),
    .Y(_0138_));
 sg13g2_nor2_1 _4586_ (.A(net677),
    .B(net729),
    .Y(_0139_));
 sg13g2_nor2_1 _4587_ (.A(net676),
    .B(net729),
    .Y(_0140_));
 sg13g2_nor2_1 _4588_ (.A(net677),
    .B(net729),
    .Y(_0141_));
 sg13g2_nor2_1 _4589_ (.A(net687),
    .B(net738),
    .Y(_0142_));
 sg13g2_nor2_1 _4590_ (.A(net687),
    .B(net738),
    .Y(_0143_));
 sg13g2_nor2_1 _4591_ (.A(net687),
    .B(net738),
    .Y(_0144_));
 sg13g2_nor2_1 _4592_ (.A(net687),
    .B(net738),
    .Y(_0145_));
 sg13g2_nor2_1 _4593_ (.A(net654),
    .B(net705),
    .Y(_0146_));
 sg13g2_nor2_1 _4594_ (.A(net655),
    .B(net706),
    .Y(_0147_));
 sg13g2_nor2_1 _4595_ (.A(net655),
    .B(net706),
    .Y(_0148_));
 sg13g2_nor2_1 _4596_ (.A(net653),
    .B(net704),
    .Y(_0149_));
 sg13g2_nor2_1 _4597_ (.A(net654),
    .B(net705),
    .Y(_0150_));
 sg13g2_nor2_1 _4598_ (.A(net653),
    .B(net704),
    .Y(_0151_));
 sg13g2_nor2_1 _4599_ (.A(net653),
    .B(net704),
    .Y(_0152_));
 sg13g2_nor2_1 _4600_ (.A(net654),
    .B(net705),
    .Y(_0153_));
 sg13g2_nor2_1 _4601_ (.A(net663),
    .B(net714),
    .Y(_0154_));
 sg13g2_nor2_1 _4602_ (.A(net666),
    .B(net717),
    .Y(_0155_));
 sg13g2_nor2_1 _4603_ (.A(net668),
    .B(net720),
    .Y(_0156_));
 sg13g2_nor2_1 _4604_ (.A(net666),
    .B(net717),
    .Y(_0157_));
 sg13g2_nor2_1 _4605_ (.A(net691),
    .B(net743),
    .Y(_0158_));
 sg13g2_nor2_1 _4606_ (.A(net691),
    .B(net743),
    .Y(_0159_));
 sg13g2_nor2_1 _4607_ (.A(net691),
    .B(net743),
    .Y(_0160_));
 sg13g2_nor2_1 _4608_ (.A(net691),
    .B(net743),
    .Y(_0161_));
 sg13g2_nor2_1 _4609_ (.A(net690),
    .B(net744),
    .Y(_0162_));
 sg13g2_nor2_1 _4610_ (.A(net690),
    .B(net744),
    .Y(_0163_));
 sg13g2_nor2_1 _4611_ (.A(net691),
    .B(net743),
    .Y(_0164_));
 sg13g2_nor2_1 _4612_ (.A(net692),
    .B(net744),
    .Y(_0165_));
 sg13g2_nor2_1 _4613_ (.A(net690),
    .B(net744),
    .Y(_0166_));
 sg13g2_nor2_1 _4614_ (.A(net691),
    .B(net743),
    .Y(_0167_));
 sg13g2_nor2_1 _4615_ (.A(net690),
    .B(net743),
    .Y(_0168_));
 sg13g2_nor2_1 _4616_ (.A(net690),
    .B(net744),
    .Y(_0169_));
 sg13g2_nor2_1 _4617_ (.A(net689),
    .B(net741),
    .Y(_0170_));
 sg13g2_nor2_1 _4618_ (.A(net689),
    .B(net741),
    .Y(_0171_));
 sg13g2_nor2_1 _4619_ (.A(net689),
    .B(net741),
    .Y(_0172_));
 sg13g2_nor2_1 _4620_ (.A(net692),
    .B(net741),
    .Y(_0173_));
 sg13g2_nor2_1 _4621_ (.A(net688),
    .B(net742),
    .Y(_0174_));
 sg13g2_nor2_1 _4622_ (.A(net688),
    .B(net740),
    .Y(_0175_));
 sg13g2_nor2_1 _4623_ (.A(net689),
    .B(net742),
    .Y(_0176_));
 sg13g2_nor2_1 _4624_ (.A(net688),
    .B(net740),
    .Y(_0177_));
 sg13g2_nor2_1 _4625_ (.A(net689),
    .B(net741),
    .Y(_0178_));
 sg13g2_nor2_1 _4626_ (.A(net688),
    .B(net740),
    .Y(_0179_));
 sg13g2_nor2_1 _4627_ (.A(net688),
    .B(net740),
    .Y(_0180_));
 sg13g2_nor2_1 _4628_ (.A(net688),
    .B(net740),
    .Y(_0181_));
 sg13g2_nor2_1 _4629_ (.A(net689),
    .B(net741),
    .Y(_0182_));
 sg13g2_nor2_1 _4630_ (.A(net692),
    .B(net740),
    .Y(_0183_));
 sg13g2_nor2_1 _4631_ (.A(net688),
    .B(net740),
    .Y(_0184_));
 sg13g2_nor2_1 _4632_ (.A(net688),
    .B(net740),
    .Y(_0185_));
 sg13g2_nor2_1 _4633_ (.A(net670),
    .B(net721),
    .Y(_0186_));
 sg13g2_nor2_1 _4634_ (.A(net670),
    .B(net721),
    .Y(_0187_));
 sg13g2_nor2_1 _4635_ (.A(net666),
    .B(net717),
    .Y(_0188_));
 sg13g2_nor2_1 _4636_ (.A(net666),
    .B(net717),
    .Y(_0189_));
 sg13g2_nor2_1 _4637_ (.A(net667),
    .B(net717),
    .Y(_0190_));
 sg13g2_nor2_1 _4638_ (.A(net666),
    .B(net717),
    .Y(_0191_));
 sg13g2_nor2_1 _4639_ (.A(net667),
    .B(net718),
    .Y(_0192_));
 sg13g2_nor2_1 _4640_ (.A(net666),
    .B(net718),
    .Y(_0193_));
 sg13g2_nor2_1 _4641_ (.A(net661),
    .B(net712),
    .Y(_0194_));
 sg13g2_nor2_1 _4642_ (.A(net664),
    .B(net715),
    .Y(_0195_));
 sg13g2_nor2_1 _4643_ (.A(net663),
    .B(net714),
    .Y(_0196_));
 sg13g2_nor2_1 _4644_ (.A(net664),
    .B(net715),
    .Y(_0197_));
 sg13g2_nor2_1 _4645_ (.A(net672),
    .B(net723),
    .Y(_0198_));
 sg13g2_nor2_1 _4646_ (.A(net670),
    .B(net721),
    .Y(_0199_));
 sg13g2_nor2_1 _4647_ (.A(net668),
    .B(net720),
    .Y(_0200_));
 sg13g2_nor2_1 _4648_ (.A(net670),
    .B(net721),
    .Y(_0201_));
 sg13g2_nor2_1 _4649_ (.A(net659),
    .B(net710),
    .Y(_0202_));
 sg13g2_nor2_1 _4650_ (.A(net668),
    .B(net719),
    .Y(_0203_));
 sg13g2_nor2_1 _4651_ (.A(net669),
    .B(net719),
    .Y(_0204_));
 sg13g2_nor2_1 _4652_ (.A(net684),
    .B(net735),
    .Y(_0205_));
 sg13g2_nor2_1 _4653_ (.A(net669),
    .B(net720),
    .Y(_0206_));
 sg13g2_nor2_1 _4654_ (.A(net684),
    .B(net719),
    .Y(_0207_));
 sg13g2_nor2_1 _4655_ (.A(net669),
    .B(net719),
    .Y(_0208_));
 sg13g2_nor2_1 _4656_ (.A(net669),
    .B(net719),
    .Y(_0209_));
 sg13g2_nor2_1 _4657_ (.A(net669),
    .B(net719),
    .Y(_0210_));
 sg13g2_nor2_1 _4658_ (.A(net684),
    .B(net719),
    .Y(_0211_));
 sg13g2_nor2_1 _4659_ (.A(net669),
    .B(net719),
    .Y(_0212_));
 sg13g2_nor2_1 _4660_ (.A(net684),
    .B(net735),
    .Y(_0213_));
 sg13g2_nor2_1 _4661_ (.A(net659),
    .B(net710),
    .Y(_0214_));
 sg13g2_nor2_1 _4662_ (.A(net659),
    .B(net710),
    .Y(_0215_));
 sg13g2_nor2_1 _4663_ (.A(net659),
    .B(net710),
    .Y(_0216_));
 sg13g2_nor2_1 _4664_ (.A(net676),
    .B(net728),
    .Y(_0217_));
 sg13g2_nor2_1 _4665_ (.A(net686),
    .B(net737),
    .Y(_0218_));
 sg13g2_nor2_1 _4666_ (.A(net671),
    .B(net722),
    .Y(_0219_));
 sg13g2_nor2_1 _4667_ (.A(net686),
    .B(net737),
    .Y(_0220_));
 sg13g2_nor2_1 _4668_ (.A(net671),
    .B(net722),
    .Y(_0221_));
 sg13g2_nor2_1 _4669_ (.A(net687),
    .B(net738),
    .Y(_0222_));
 sg13g2_nor2_1 _4670_ (.A(net671),
    .B(net722),
    .Y(_0223_));
 sg13g2_nor2_1 _4671_ (.A(net686),
    .B(net737),
    .Y(_0224_));
 sg13g2_nor2_1 _4672_ (.A(net671),
    .B(net722),
    .Y(_0225_));
 sg13g2_nor2_1 _4673_ (.A(net686),
    .B(net738),
    .Y(_0226_));
 sg13g2_nor2_1 _4674_ (.A(net671),
    .B(net723),
    .Y(_0227_));
 sg13g2_nor2_1 _4675_ (.A(net686),
    .B(net737),
    .Y(_0228_));
 sg13g2_nor2_1 _4676_ (.A(net671),
    .B(net722),
    .Y(_0229_));
 sg13g2_nor2_1 _4677_ (.A(net671),
    .B(net722),
    .Y(_0230_));
 sg13g2_nor2_1 _4678_ (.A(net672),
    .B(net722),
    .Y(_0231_));
 sg13g2_nor2_1 _4679_ (.A(net686),
    .B(net737),
    .Y(_0232_));
 sg13g2_nor2_1 _4680_ (.A(net671),
    .B(net722),
    .Y(_0233_));
 sg13g2_nor2_1 _4681_ (.A(net663),
    .B(net714),
    .Y(_0234_));
 sg13g2_nor2_1 _4682_ (.A(net664),
    .B(net715),
    .Y(_0235_));
 sg13g2_nor2_1 _4683_ (.A(net668),
    .B(net714),
    .Y(_0236_));
 sg13g2_nor2_1 _4684_ (.A(net666),
    .B(net717),
    .Y(_0237_));
 sg13g2_nor2_1 _4685_ (.A(net687),
    .B(net739),
    .Y(_0238_));
 sg13g2_nor2_1 _4686_ (.A(net685),
    .B(net735),
    .Y(_0239_));
 sg13g2_nor2_1 _4687_ (.A(net687),
    .B(net738),
    .Y(_0240_));
 sg13g2_nor2_1 _4688_ (.A(net685),
    .B(net735),
    .Y(_0241_));
 sg13g2_nor2_1 _4689_ (.A(net686),
    .B(net737),
    .Y(_0242_));
 sg13g2_nor2_1 _4690_ (.A(net685),
    .B(net736),
    .Y(_0243_));
 sg13g2_nor2_1 _4691_ (.A(net684),
    .B(net735),
    .Y(_0244_));
 sg13g2_nor2_1 _4692_ (.A(net684),
    .B(net735),
    .Y(_0245_));
 sg13g2_nor2_1 _4693_ (.A(net661),
    .B(net712),
    .Y(_0246_));
 sg13g2_nor2_1 _4694_ (.A(net665),
    .B(net716),
    .Y(_0247_));
 sg13g2_nor2_1 _4695_ (.A(net662),
    .B(net713),
    .Y(_0248_));
 sg13g2_nor2_1 _4696_ (.A(net664),
    .B(net715),
    .Y(_0249_));
 sg13g2_nor2_1 _4697_ (.A(net690),
    .B(net744),
    .Y(_0250_));
 sg13g2_nor2_1 _4698_ (.A(net690),
    .B(net744),
    .Y(_0251_));
 sg13g2_nor2_1 _4699_ (.A(net691),
    .B(net743),
    .Y(_0252_));
 sg13g2_nor2_1 _4700_ (.A(net690),
    .B(net744),
    .Y(_0253_));
 sg13g2_nor2_1 _4701_ (.A(net661),
    .B(net712),
    .Y(_0254_));
 sg13g2_nor2_1 _4702_ (.A(net665),
    .B(net716),
    .Y(_0255_));
 sg13g2_nor2_1 _4703_ (.A(net662),
    .B(net713),
    .Y(_0256_));
 sg13g2_nor2_1 _4704_ (.A(net665),
    .B(net716),
    .Y(_0257_));
 sg13g2_nor2_1 _4705_ (.A(_1994_),
    .B(_1998_),
    .Y(_0613_));
 sg13g2_nor2_1 _4706_ (.A(_1994_),
    .B(_1998_),
    .Y(_0614_));
 sg13g2_nor2_1 _4707_ (.A(net654),
    .B(net705),
    .Y(_0258_));
 sg13g2_nor2_1 _4708_ (.A(net653),
    .B(net704),
    .Y(_0259_));
 sg13g2_nor2_1 _4709_ (.A(net656),
    .B(net707),
    .Y(_0260_));
 sg13g2_nor2_1 _4710_ (.A(net653),
    .B(net704),
    .Y(_0261_));
 sg13g2_dfrbpq_1 _4711_ (.RESET_B(net253),
    .D(_0263_),
    .Q(\tmds_green.dc_balancing_reg[0] ),
    .CLK(net648));
 sg13g2_dfrbpq_1 _4712_ (.RESET_B(net156),
    .D(_0264_),
    .Q(\tmds_blue.dc_balancing_reg[0] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4713_ (.RESET_B(net154),
    .D(_0265_),
    .Q(\clockdiv.q1 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _4714_ (.RESET_B(net153),
    .D(_0266_),
    .Q(\clockdiv.q2 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _4715_ (.RESET_B(net152),
    .D(net737),
    .Q(\clockdiv.q2temp ),
    .CLK(net405));
 sg13g2_dfrbpq_1 _4716_ (.RESET_B(net151),
    .D(_0267_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ),
    .CLK(_0006_));
 sg13g2_dfrbpq_1 _4717_ (.RESET_B(net149),
    .D(_0268_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .CLK(_0007_));
 sg13g2_dfrbpq_1 _4718_ (.RESET_B(net147),
    .D(_0269_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .CLK(_0008_));
 sg13g2_dfrbpq_1 _4719_ (.RESET_B(net145),
    .D(_0270_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .CLK(_0009_));
 sg13g2_dfrbpq_1 _4720_ (.RESET_B(net143),
    .D(_0271_),
    .Q(\green_tmds_par[0] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _4721_ (.RESET_B(net142),
    .D(_0272_),
    .Q(\green_tmds_par[1] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _4722_ (.RESET_B(net141),
    .D(_0273_),
    .Q(\green_tmds_par[7] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _4723_ (.RESET_B(net140),
    .D(_0274_),
    .Q(\red_tmds_par[0] ),
    .CLK(net647));
 sg13g2_dfrbpq_1 _4724_ (.RESET_B(net139),
    .D(_0275_),
    .Q(\red_tmds_par[1] ),
    .CLK(net647));
 sg13g2_dfrbpq_1 _4725_ (.RESET_B(net138),
    .D(_0276_),
    .Q(\red_tmds_par[3] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4726_ (.RESET_B(net137),
    .D(_0277_),
    .Q(\red_tmds_par[5] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4727_ (.RESET_B(net136),
    .D(_0278_),
    .Q(\red_tmds_par[7] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4728_ (.RESET_B(net135),
    .D(_0279_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .CLK(_0010_));
 sg13g2_dfrbpq_1 _4729_ (.RESET_B(net133),
    .D(_0280_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ),
    .CLK(_0011_));
 sg13g2_dfrbpq_1 _4730_ (.RESET_B(net131),
    .D(_0281_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .CLK(_0012_));
 sg13g2_dfrbpq_1 _4731_ (.RESET_B(net129),
    .D(_0282_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ),
    .CLK(_0013_));
 sg13g2_dfrbpq_1 _4732_ (.RESET_B(net127),
    .D(_0283_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .CLK(_0014_));
 sg13g2_dfrbpq_1 _4733_ (.RESET_B(net125),
    .D(_0284_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .CLK(_0015_));
 sg13g2_dfrbpq_1 _4734_ (.RESET_B(net123),
    .D(_0285_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .CLK(_0016_));
 sg13g2_dfrbpq_1 _4735_ (.RESET_B(net121),
    .D(_0286_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .CLK(_0017_));
 sg13g2_dfrbpq_1 _4736_ (.RESET_B(net119),
    .D(_0287_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .CLK(_0018_));
 sg13g2_dfrbpq_1 _4737_ (.RESET_B(net117),
    .D(_0288_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .CLK(_0019_));
 sg13g2_dfrbpq_1 _4738_ (.RESET_B(net115),
    .D(_0289_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .CLK(_0020_));
 sg13g2_dfrbpq_1 _4739_ (.RESET_B(net113),
    .D(_0290_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .CLK(_0021_));
 sg13g2_dfrbpq_1 _4740_ (.RESET_B(net111),
    .D(_0291_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .CLK(_0022_));
 sg13g2_dfrbpq_1 _4741_ (.RESET_B(net109),
    .D(_0292_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .CLK(_0023_));
 sg13g2_dfrbpq_1 _4742_ (.RESET_B(net107),
    .D(_0293_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .CLK(_0024_));
 sg13g2_dfrbpq_1 _4743_ (.RESET_B(net105),
    .D(_0294_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .CLK(_0025_));
 sg13g2_dfrbpq_1 _4744_ (.RESET_B(net103),
    .D(_0295_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .CLK(_0026_));
 sg13g2_dfrbpq_1 _4745_ (.RESET_B(net101),
    .D(_0296_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .CLK(_0027_));
 sg13g2_dfrbpq_1 _4746_ (.RESET_B(net99),
    .D(_0297_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .CLK(_0028_));
 sg13g2_dfrbpq_1 _4747_ (.RESET_B(net97),
    .D(_0298_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .CLK(_0029_));
 sg13g2_dfrbpq_1 _4748_ (.RESET_B(net95),
    .D(_0299_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .CLK(_0030_));
 sg13g2_dfrbpq_1 _4749_ (.RESET_B(net93),
    .D(_0300_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .CLK(_0031_));
 sg13g2_dfrbpq_1 _4750_ (.RESET_B(net91),
    .D(_0301_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .CLK(_0032_));
 sg13g2_dfrbpq_1 _4751_ (.RESET_B(net89),
    .D(_0302_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .CLK(_0033_));
 sg13g2_dfrbpq_2 _4752_ (.RESET_B(net87),
    .D(_0303_),
    .Q(\videogen.fancy_shader.video_x[0] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4753_ (.RESET_B(net86),
    .D(_0304_),
    .Q(\videogen.fancy_shader.video_x[1] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4754_ (.RESET_B(net85),
    .D(_0305_),
    .Q(\videogen.fancy_shader.video_x[2] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _4755_ (.RESET_B(net84),
    .D(_0306_),
    .Q(\videogen.fancy_shader.video_x[3] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _4756_ (.RESET_B(net83),
    .D(_0307_),
    .Q(\videogen.fancy_shader.video_x[4] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4757_ (.RESET_B(net82),
    .D(_0308_),
    .Q(\videogen.fancy_shader.video_x[5] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4758_ (.RESET_B(net81),
    .D(_0309_),
    .Q(\videogen.fancy_shader.video_x[6] ),
    .CLK(net638));
 sg13g2_dfrbpq_1 _4759_ (.RESET_B(net80),
    .D(_0310_),
    .Q(\videogen.fancy_shader.video_x[7] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4760_ (.RESET_B(net79),
    .D(_0311_),
    .Q(\videogen.fancy_shader.video_x[8] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4761_ (.RESET_B(net78),
    .D(_0312_),
    .Q(\videogen.fancy_shader.video_x[9] ),
    .CLK(net638));
 sg13g2_dfrbpq_1 _4762_ (.RESET_B(net77),
    .D(_0313_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .CLK(_0034_));
 sg13g2_dfrbpq_1 _4763_ (.RESET_B(net75),
    .D(_0314_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .CLK(_0035_));
 sg13g2_dfrbpq_1 _4764_ (.RESET_B(net73),
    .D(_0315_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .CLK(_0036_));
 sg13g2_dfrbpq_1 _4765_ (.RESET_B(net71),
    .D(_0316_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .CLK(_0037_));
 sg13g2_dfrbpq_1 _4766_ (.RESET_B(net69),
    .D(_0317_),
    .Q(\tmds_blue.vsync ),
    .CLK(net640));
 sg13g2_dfrbpq_2 _4767_ (.RESET_B(net68),
    .D(_0318_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4768_ (.RESET_B(net66),
    .D(_0319_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4769_ (.RESET_B(net64),
    .D(_0320_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4770_ (.RESET_B(net62),
    .D(_0321_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4771_ (.RESET_B(net60),
    .D(_0322_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4772_ (.RESET_B(net58),
    .D(_0323_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4773_ (.RESET_B(net56),
    .D(_0324_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ),
    .CLK(net633));
 sg13g2_dfrbpq_1 _4774_ (.RESET_B(net54),
    .D(_0325_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .CLK(net633));
 sg13g2_dfrbpq_1 _4775_ (.RESET_B(net52),
    .D(_0326_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4776_ (.RESET_B(net50),
    .D(_0327_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4777_ (.RESET_B(net48),
    .D(_0328_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4778_ (.RESET_B(net46),
    .D(_0329_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .CLK(net632));
 sg13g2_dfrbpq_1 _4779_ (.RESET_B(net44),
    .D(_0330_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4780_ (.RESET_B(net42),
    .D(_0331_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4781_ (.RESET_B(net40),
    .D(_0332_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4782_ (.RESET_B(net38),
    .D(_0333_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .CLK(net632));
 sg13g2_dfrbpq_1 _4783_ (.RESET_B(net36),
    .D(_0334_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .CLK(net633));
 sg13g2_dfrbpq_1 _4784_ (.RESET_B(net34),
    .D(_0335_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4785_ (.RESET_B(net32),
    .D(_0336_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .CLK(net633));
 sg13g2_dfrbpq_1 _4786_ (.RESET_B(net404),
    .D(_0337_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4787_ (.RESET_B(net400),
    .D(_0338_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .CLK(_0038_));
 sg13g2_dfrbpq_1 _4788_ (.RESET_B(net398),
    .D(_0339_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .CLK(_0039_));
 sg13g2_dfrbpq_1 _4789_ (.RESET_B(net396),
    .D(_0340_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .CLK(_0040_));
 sg13g2_dfrbpq_1 _4790_ (.RESET_B(net394),
    .D(_0341_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .CLK(_0041_));
 sg13g2_dfrbpq_1 _4791_ (.RESET_B(net392),
    .D(_0342_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .CLK(_0042_));
 sg13g2_dfrbpq_1 _4792_ (.RESET_B(net390),
    .D(_0343_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .CLK(_0043_));
 sg13g2_dfrbpq_1 _4793_ (.RESET_B(net388),
    .D(_0344_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .CLK(_0044_));
 sg13g2_dfrbpq_1 _4794_ (.RESET_B(net386),
    .D(_0345_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .CLK(_0045_));
 sg13g2_dfrbpq_2 _4795_ (.RESET_B(net384),
    .D(_0346_),
    .Q(\videogen.fancy_shader.n646[0] ),
    .CLK(net649));
 sg13g2_dfrbpq_2 _4796_ (.RESET_B(net382),
    .D(_0347_),
    .Q(\videogen.fancy_shader.n646[1] ),
    .CLK(net649));
 sg13g2_dfrbpq_2 _4797_ (.RESET_B(net380),
    .D(_0348_),
    .Q(\videogen.fancy_shader.n646[2] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _4798_ (.RESET_B(net378),
    .D(_0349_),
    .Q(\videogen.fancy_shader.n646[3] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4799_ (.RESET_B(net376),
    .D(_0350_),
    .Q(\videogen.fancy_shader.n646[4] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _4800_ (.RESET_B(net374),
    .D(_0351_),
    .Q(\videogen.fancy_shader.n646[5] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4801_ (.RESET_B(net372),
    .D(_0352_),
    .Q(\videogen.fancy_shader.n646[6] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _4802_ (.RESET_B(net370),
    .D(_0353_),
    .Q(\videogen.fancy_shader.n646[7] ),
    .CLK(net633));
 sg13g2_dfrbpq_1 _4803_ (.RESET_B(net368),
    .D(_0354_),
    .Q(\videogen.fancy_shader.n646[8] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4804_ (.RESET_B(net366),
    .D(_0355_),
    .Q(\videogen.fancy_shader.n646[9] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4805_ (.RESET_B(net364),
    .D(_0356_),
    .Q(\videogen.fancy_shader.video_y[0] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _4806_ (.RESET_B(net362),
    .D(_0357_),
    .Q(\videogen.fancy_shader.video_y[1] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _4807_ (.RESET_B(net360),
    .D(_0358_),
    .Q(\videogen.fancy_shader.video_y[2] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4808_ (.RESET_B(net358),
    .D(_0359_),
    .Q(\videogen.fancy_shader.video_y[3] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4809_ (.RESET_B(net356),
    .D(_0360_),
    .Q(\videogen.fancy_shader.video_y[4] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4810_ (.RESET_B(net354),
    .D(_0361_),
    .Q(\videogen.fancy_shader.video_y[5] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4811_ (.RESET_B(net352),
    .D(_0362_),
    .Q(\videogen.fancy_shader.video_y[6] ),
    .CLK(net635));
 sg13g2_dfrbpq_2 _4812_ (.RESET_B(net350),
    .D(_0363_),
    .Q(\videogen.fancy_shader.video_y[7] ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4813_ (.RESET_B(net348),
    .D(_0364_),
    .Q(\videogen.fancy_shader.video_y[8] ),
    .CLK(net635));
 sg13g2_dfrbpq_2 _4814_ (.RESET_B(net346),
    .D(_0365_),
    .Q(\videogen.fancy_shader.video_y[9] ),
    .CLK(net635));
 sg13g2_dfrbpq_2 _4815_ (.RESET_B(net344),
    .D(_0366_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .CLK(net643));
 sg13g2_dfrbpq_2 _4816_ (.RESET_B(net343),
    .D(_0367_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _4817_ (.RESET_B(net342),
    .D(_0368_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[2] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _4818_ (.RESET_B(net341),
    .D(_0369_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .CLK(net643));
 sg13g2_dfrbpq_2 _4819_ (.RESET_B(net340),
    .D(_0370_),
    .Q(hsync),
    .CLK(net640));
 sg13g2_dfrbpq_1 _4820_ (.RESET_B(net339),
    .D(_0371_),
    .Q(display_enable),
    .CLK(net640));
 sg13g2_dfrbpq_2 _4821_ (.RESET_B(net338),
    .D(_0372_),
    .Q(\tmds_blue.n193 ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4822_ (.RESET_B(net337),
    .D(_0373_),
    .Q(\tmds_blue.n100 ),
    .CLK(net640));
 sg13g2_dfrbpq_1 _4823_ (.RESET_B(net336),
    .D(_0374_),
    .Q(\tmds_blue.n126 ),
    .CLK(net640));
 sg13g2_dfrbpq_2 _4824_ (.RESET_B(net335),
    .D(_0375_),
    .Q(\tmds_blue.n132 ),
    .CLK(net640));
 sg13g2_dfrbpq_2 _4825_ (.RESET_B(net334),
    .D(_0376_),
    .Q(\tmds_green.n100 ),
    .CLK(net642));
 sg13g2_dfrbpq_2 _4826_ (.RESET_B(net333),
    .D(_0377_),
    .Q(\tmds_green.n126 ),
    .CLK(net640));
 sg13g2_dfrbpq_1 _4827_ (.RESET_B(net332),
    .D(_0378_),
    .Q(\tmds_green.n132 ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4828_ (.RESET_B(net331),
    .D(_0379_),
    .Q(\tmds_red.n102 ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _4829_ (.RESET_B(net330),
    .D(_0380_),
    .Q(\tmds_red.n100 ),
    .CLK(net649));
 sg13g2_dfrbpq_2 _4830_ (.RESET_B(net329),
    .D(_0381_),
    .Q(\tmds_red.n114 ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _4831_ (.RESET_B(net328),
    .D(_0382_),
    .Q(\tmds_red.n126 ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _4832_ (.RESET_B(net327),
    .D(_0383_),
    .Q(\tmds_red.n132 ),
    .CLK(net640));
 sg13g2_dfrbpq_1 _4833_ (.RESET_B(net326),
    .D(_0384_),
    .Q(\red_tmds_par[2] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4834_ (.RESET_B(net325),
    .D(_0385_),
    .Q(\red_tmds_par[4] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4835_ (.RESET_B(net324),
    .D(_0386_),
    .Q(\red_tmds_par[6] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4836_ (.RESET_B(net323),
    .D(_0387_),
    .Q(\red_tmds_par[8] ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _4837_ (.RESET_B(net322),
    .D(_0388_),
    .Q(\red_tmds_par[9] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4838_ (.RESET_B(net321),
    .D(_0389_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .CLK(_0046_));
 sg13g2_dfrbpq_1 _4839_ (.RESET_B(net319),
    .D(_0390_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .CLK(_0047_));
 sg13g2_dfrbpq_1 _4840_ (.RESET_B(net317),
    .D(_0391_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .CLK(_0048_));
 sg13g2_dfrbpq_1 _4841_ (.RESET_B(net315),
    .D(_0392_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .CLK(_0049_));
 sg13g2_dfrbpq_1 _4842_ (.RESET_B(net313),
    .D(_0393_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .CLK(_0050_));
 sg13g2_dfrbpq_1 _4843_ (.RESET_B(net311),
    .D(_0394_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .CLK(_0051_));
 sg13g2_dfrbpq_1 _4844_ (.RESET_B(net309),
    .D(_0395_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .CLK(_0052_));
 sg13g2_dfrbpq_1 _4845_ (.RESET_B(net307),
    .D(_0396_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .CLK(_0053_));
 sg13g2_dfrbpq_1 _4846_ (.RESET_B(net305),
    .D(_0397_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ),
    .CLK(_0054_));
 sg13g2_dfrbpq_1 _4847_ (.RESET_B(net303),
    .D(_0398_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ),
    .CLK(_0055_));
 sg13g2_dfrbpq_1 _4848_ (.RESET_B(net301),
    .D(_0399_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ),
    .CLK(_0056_));
 sg13g2_dfrbpq_1 _4849_ (.RESET_B(net299),
    .D(_0400_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .CLK(_0057_));
 sg13g2_dfrbpq_1 _4850_ (.RESET_B(net298),
    .D(_0401_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .CLK(_0058_));
 sg13g2_dfrbpq_1 _4851_ (.RESET_B(net296),
    .D(_0402_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .CLK(_0059_));
 sg13g2_dfrbpq_1 _4852_ (.RESET_B(net294),
    .D(_0403_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .CLK(_0060_));
 sg13g2_dfrbpq_1 _4853_ (.RESET_B(net292),
    .D(_0404_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .CLK(_0061_));
 sg13g2_dfrbpq_1 _4854_ (.RESET_B(net290),
    .D(_0405_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .CLK(_0062_));
 sg13g2_dfrbpq_1 _4855_ (.RESET_B(net288),
    .D(_0406_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .CLK(_0063_));
 sg13g2_dfrbpq_1 _4856_ (.RESET_B(net286),
    .D(_0407_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .CLK(_0064_));
 sg13g2_dfrbpq_1 _4857_ (.RESET_B(net284),
    .D(_0408_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .CLK(_0065_));
 sg13g2_dfrbpq_1 _4858_ (.RESET_B(net282),
    .D(_0409_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .CLK(_0066_));
 sg13g2_dfrbpq_1 _4859_ (.RESET_B(net280),
    .D(_0410_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ),
    .CLK(_0067_));
 sg13g2_dfrbpq_1 _4860_ (.RESET_B(net278),
    .D(_0411_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .CLK(_0068_));
 sg13g2_dfrbpq_1 _4861_ (.RESET_B(net276),
    .D(_0412_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .CLK(_0069_));
 sg13g2_dfrbpq_1 _4862_ (.RESET_B(net274),
    .D(_0413_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ),
    .CLK(_0070_));
 sg13g2_dfrbpq_1 _4863_ (.RESET_B(net272),
    .D(_0414_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .CLK(_0071_));
 sg13g2_dfrbpq_1 _4864_ (.RESET_B(net270),
    .D(_0415_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .CLK(_0072_));
 sg13g2_dfrbpq_1 _4865_ (.RESET_B(net268),
    .D(_0416_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .CLK(_0073_));
 sg13g2_dfrbpq_1 _4866_ (.RESET_B(net267),
    .D(_0417_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ),
    .CLK(_0074_));
 sg13g2_dfrbpq_1 _4867_ (.RESET_B(net265),
    .D(_0418_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .CLK(_0075_));
 sg13g2_dfrbpq_1 _4868_ (.RESET_B(net263),
    .D(_0419_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .CLK(_0076_));
 sg13g2_dfrbpq_1 _4869_ (.RESET_B(net261),
    .D(_0420_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .CLK(_0077_));
 sg13g2_dfrbpq_1 _4870_ (.RESET_B(net259),
    .D(_0421_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .CLK(_0078_));
 sg13g2_dfrbpq_1 _4871_ (.RESET_B(net257),
    .D(_0422_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .CLK(_0079_));
 sg13g2_dfrbpq_1 _4872_ (.RESET_B(net251),
    .D(_0423_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .CLK(_0080_));
 sg13g2_dfrbpq_1 _4873_ (.RESET_B(net249),
    .D(_0424_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .CLK(_0081_));
 sg13g2_dfrbpq_1 _4874_ (.RESET_B(net247),
    .D(_0425_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .CLK(_0082_));
 sg13g2_dfrbpq_1 _4875_ (.RESET_B(net245),
    .D(_0426_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .CLK(_0083_));
 sg13g2_dfrbpq_1 _4876_ (.RESET_B(net243),
    .D(_0427_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .CLK(_0084_));
 sg13g2_dfrbpq_1 _4877_ (.RESET_B(net241),
    .D(_0428_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .CLK(_0085_));
 sg13g2_dfrbpq_1 _4878_ (.RESET_B(net239),
    .D(_0429_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ),
    .CLK(_0086_));
 sg13g2_dfrbpq_1 _4879_ (.RESET_B(net237),
    .D(_0430_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .CLK(_0087_));
 sg13g2_dfrbpq_1 _4880_ (.RESET_B(net235),
    .D(_0431_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .CLK(_0088_));
 sg13g2_dfrbpq_1 _4881_ (.RESET_B(net233),
    .D(_0432_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .CLK(_0089_));
 sg13g2_dfrbpq_1 _4882_ (.RESET_B(net232),
    .D(_0433_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .CLK(_0090_));
 sg13g2_dfrbpq_1 _4883_ (.RESET_B(net230),
    .D(_0434_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ),
    .CLK(_0091_));
 sg13g2_dfrbpq_1 _4884_ (.RESET_B(net228),
    .D(_0435_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .CLK(_0092_));
 sg13g2_dfrbpq_1 _4885_ (.RESET_B(net226),
    .D(_0436_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .CLK(_0093_));
 sg13g2_dfrbpq_1 _4886_ (.RESET_B(net224),
    .D(_0437_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .CLK(_0094_));
 sg13g2_dfrbpq_1 _4887_ (.RESET_B(net222),
    .D(_0438_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .CLK(_0095_));
 sg13g2_dfrbpq_1 _4888_ (.RESET_B(net220),
    .D(_0439_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .CLK(_0096_));
 sg13g2_dfrbpq_1 _4889_ (.RESET_B(net218),
    .D(_0440_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .CLK(_0097_));
 sg13g2_dfrbpq_1 _4890_ (.RESET_B(net216),
    .D(_0441_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .CLK(_0098_));
 sg13g2_dfrbpq_1 _4891_ (.RESET_B(net214),
    .D(_0442_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .CLK(_0099_));
 sg13g2_dfrbpq_1 _4892_ (.RESET_B(net212),
    .D(_0443_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .CLK(_0100_));
 sg13g2_dfrbpq_1 _4893_ (.RESET_B(net210),
    .D(_0444_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .CLK(_0101_));
 sg13g2_dfrbpq_1 _4894_ (.RESET_B(net208),
    .D(_0445_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .CLK(_0102_));
 sg13g2_dfrbpq_1 _4895_ (.RESET_B(net206),
    .D(_0446_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .CLK(_0103_));
 sg13g2_dfrbpq_1 _4896_ (.RESET_B(net204),
    .D(_0447_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .CLK(_0104_));
 sg13g2_dfrbpq_1 _4897_ (.RESET_B(net202),
    .D(_0448_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .CLK(_0105_));
 sg13g2_dfrbpq_1 _4898_ (.RESET_B(net200),
    .D(_0449_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .CLK(_0106_));
 sg13g2_dfrbpq_1 _4899_ (.RESET_B(net198),
    .D(_0450_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .CLK(_0107_));
 sg13g2_dfrbpq_1 _4900_ (.RESET_B(net196),
    .D(_0451_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .CLK(_0108_));
 sg13g2_dfrbpq_1 _4901_ (.RESET_B(net194),
    .D(_0452_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ),
    .CLK(_0109_));
 sg13g2_dfrbpq_1 _4902_ (.RESET_B(net192),
    .D(_0453_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ),
    .CLK(_0110_));
 sg13g2_dfrbpq_1 _4903_ (.RESET_B(net190),
    .D(_0454_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .CLK(_0111_));
 sg13g2_dfrbpq_1 _4904_ (.RESET_B(net188),
    .D(_0455_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .CLK(_0112_));
 sg13g2_dfrbpq_1 _4905_ (.RESET_B(net186),
    .D(_0456_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .CLK(_0113_));
 sg13g2_dfrbpq_1 _4906_ (.RESET_B(net184),
    .D(_0457_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ),
    .CLK(_0114_));
 sg13g2_dfrbpq_1 _4907_ (.RESET_B(net182),
    .D(_0458_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .CLK(_0115_));
 sg13g2_dfrbpq_1 _4908_ (.RESET_B(net180),
    .D(_0459_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .CLK(_0116_));
 sg13g2_dfrbpq_1 _4909_ (.RESET_B(net178),
    .D(_0460_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .CLK(_0117_));
 sg13g2_dfrbpq_1 _4910_ (.RESET_B(net176),
    .D(_0461_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .CLK(_0118_));
 sg13g2_dfrbpq_1 _4911_ (.RESET_B(net174),
    .D(_0462_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .CLK(_0119_));
 sg13g2_dfrbpq_1 _4912_ (.RESET_B(net172),
    .D(_0463_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .CLK(_0120_));
 sg13g2_dfrbpq_1 _4913_ (.RESET_B(net170),
    .D(_0464_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ),
    .CLK(_0121_));
 sg13g2_dfrbpq_1 _4914_ (.RESET_B(net168),
    .D(_0465_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .CLK(_0122_));
 sg13g2_dfrbpq_1 _4915_ (.RESET_B(net166),
    .D(_0466_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .CLK(_0123_));
 sg13g2_dfrbpq_1 _4916_ (.RESET_B(net164),
    .D(_0467_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .CLK(_0124_));
 sg13g2_dfrbpq_1 _4917_ (.RESET_B(net162),
    .D(_0468_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .CLK(_0125_));
 sg13g2_dfrbpq_1 _4918_ (.RESET_B(net160),
    .D(_0469_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .CLK(_0126_));
 sg13g2_dfrbpq_1 _4919_ (.RESET_B(net158),
    .D(_0470_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .CLK(_0127_));
 sg13g2_dfrbpq_1 _4920_ (.RESET_B(net155),
    .D(_0471_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .CLK(_0128_));
 sg13g2_dfrbpq_1 _4921_ (.RESET_B(net148),
    .D(_0472_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .CLK(_0129_));
 sg13g2_dfrbpq_1 _4922_ (.RESET_B(net144),
    .D(_0473_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ),
    .CLK(_0130_));
 sg13g2_dfrbpq_1 _4923_ (.RESET_B(net132),
    .D(_0474_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ),
    .CLK(_0131_));
 sg13g2_dfrbpq_1 _4924_ (.RESET_B(net128),
    .D(_0475_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .CLK(_0132_));
 sg13g2_dfrbpq_1 _4925_ (.RESET_B(net124),
    .D(_0476_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .CLK(_0133_));
 sg13g2_dfrbpq_1 _4926_ (.RESET_B(net120),
    .D(_0477_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .CLK(_0134_));
 sg13g2_dfrbpq_1 _4927_ (.RESET_B(net116),
    .D(_0478_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .CLK(_0135_));
 sg13g2_dfrbpq_1 _4928_ (.RESET_B(net112),
    .D(_0479_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .CLK(_0136_));
 sg13g2_dfrbpq_1 _4929_ (.RESET_B(net108),
    .D(_0480_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .CLK(_0137_));
 sg13g2_dfrbpq_1 _4930_ (.RESET_B(net104),
    .D(_0481_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ),
    .CLK(_0138_));
 sg13g2_dfrbpq_1 _4931_ (.RESET_B(net100),
    .D(_0482_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ),
    .CLK(_0139_));
 sg13g2_dfrbpq_1 _4932_ (.RESET_B(net96),
    .D(_0483_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .CLK(_0140_));
 sg13g2_dfrbpq_1 _4933_ (.RESET_B(net254),
    .D(_0484_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .CLK(_0141_));
 sg13g2_dfrbpq_1 _4934_ (.RESET_B(net255),
    .D(_0002_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _4935_ (.RESET_B(net256),
    .D(_0003_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4936_ (.RESET_B(net402),
    .D(_0000_),
    .Q(\videogen.mem_read ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4937_ (.RESET_B(net92),
    .D(_0001_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[3] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4938_ (.RESET_B(net88),
    .D(_0485_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ),
    .CLK(_0142_));
 sg13g2_dfrbpq_1 _4939_ (.RESET_B(net74),
    .D(_0486_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ),
    .CLK(_0143_));
 sg13g2_dfrbpq_1 _4940_ (.RESET_B(net70),
    .D(_0487_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .CLK(_0144_));
 sg13g2_dfrbpq_1 _4941_ (.RESET_B(net65),
    .D(_0488_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ),
    .CLK(_0145_));
 sg13g2_dfrbpq_1 _4942_ (.RESET_B(net61),
    .D(_0489_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .CLK(_0146_));
 sg13g2_dfrbpq_1 _4943_ (.RESET_B(net57),
    .D(_0490_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .CLK(_0147_));
 sg13g2_dfrbpq_1 _4944_ (.RESET_B(net53),
    .D(_0491_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .CLK(_0148_));
 sg13g2_dfrbpq_1 _4945_ (.RESET_B(net49),
    .D(_0492_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .CLK(_0149_));
 sg13g2_dfrbpq_1 _4946_ (.RESET_B(net45),
    .D(_0493_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .CLK(_0150_));
 sg13g2_dfrbpq_1 _4947_ (.RESET_B(net41),
    .D(_0494_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .CLK(_0151_));
 sg13g2_dfrbpq_1 _4948_ (.RESET_B(net37),
    .D(_0495_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .CLK(_0152_));
 sg13g2_dfrbpq_1 _4949_ (.RESET_B(net33),
    .D(_0496_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .CLK(_0153_));
 sg13g2_dfrbpq_1 _4950_ (.RESET_B(net401),
    .D(_0497_),
    .Q(\green_tmds_par[2] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4951_ (.RESET_B(net399),
    .D(_0498_),
    .Q(\green_tmds_par[6] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4952_ (.RESET_B(net397),
    .D(_0499_),
    .Q(\green_tmds_par[8] ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _4953_ (.RESET_B(net395),
    .D(_0500_),
    .Q(\green_tmds_par[9] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _4954_ (.RESET_B(net393),
    .D(_0501_),
    .Q(\tmds_red.dc_balancing_reg[0] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4955_ (.RESET_B(net391),
    .D(_0502_),
    .Q(\tmds_red.dc_balancing_reg[1] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4956_ (.RESET_B(net389),
    .D(_0503_),
    .Q(\tmds_red.dc_balancing_reg[2] ),
    .CLK(net647));
 sg13g2_dfrbpq_1 _4957_ (.RESET_B(net387),
    .D(_0504_),
    .Q(\tmds_red.dc_balancing_reg[3] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4958_ (.RESET_B(net385),
    .D(_0505_),
    .Q(\tmds_red.dc_balancing_reg[4] ),
    .CLK(net647));
 sg13g2_dfrbpq_1 _4959_ (.RESET_B(net383),
    .D(_0506_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .CLK(_0154_));
 sg13g2_dfrbpq_1 _4960_ (.RESET_B(net379),
    .D(_0507_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .CLK(_0155_));
 sg13g2_dfrbpq_1 _4961_ (.RESET_B(net375),
    .D(_0508_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .CLK(_0156_));
 sg13g2_dfrbpq_1 _4962_ (.RESET_B(net371),
    .D(_0509_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ),
    .CLK(_0157_));
 sg13g2_dfrbpq_1 _4963_ (.RESET_B(net367),
    .D(_0510_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .CLK(_0158_));
 sg13g2_dfrbpq_1 _4964_ (.RESET_B(net363),
    .D(_0511_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .CLK(_0159_));
 sg13g2_dfrbpq_1 _4965_ (.RESET_B(net359),
    .D(_0512_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .CLK(_0160_));
 sg13g2_dfrbpq_1 _4966_ (.RESET_B(net355),
    .D(_0513_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .CLK(_0161_));
 sg13g2_dfrbpq_1 _4967_ (.RESET_B(net351),
    .D(_0514_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .CLK(_0162_));
 sg13g2_dfrbpq_1 _4968_ (.RESET_B(net347),
    .D(_0515_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .CLK(_0163_));
 sg13g2_dfrbpq_1 _4969_ (.RESET_B(net320),
    .D(_0516_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .CLK(_0164_));
 sg13g2_dfrbpq_1 _4970_ (.RESET_B(net316),
    .D(_0517_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .CLK(_0165_));
 sg13g2_dfrbpq_1 _4971_ (.RESET_B(net312),
    .D(_0518_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .CLK(_0166_));
 sg13g2_dfrbpq_1 _4972_ (.RESET_B(net308),
    .D(_0519_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .CLK(_0167_));
 sg13g2_dfrbpq_1 _4973_ (.RESET_B(net304),
    .D(_0520_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .CLK(_0168_));
 sg13g2_dfrbpq_1 _4974_ (.RESET_B(net300),
    .D(_0521_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .CLK(_0169_));
 sg13g2_dfrbpq_1 _4975_ (.RESET_B(net297),
    .D(_0522_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ),
    .CLK(_0170_));
 sg13g2_dfrbpq_1 _4976_ (.RESET_B(net293),
    .D(_0523_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ),
    .CLK(_0171_));
 sg13g2_dfrbpq_1 _4977_ (.RESET_B(net289),
    .D(_0524_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .CLK(_0172_));
 sg13g2_dfrbpq_1 _4978_ (.RESET_B(net285),
    .D(_0525_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .CLK(_0173_));
 sg13g2_dfrbpq_1 _4979_ (.RESET_B(net281),
    .D(_0526_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .CLK(_0174_));
 sg13g2_dfrbpq_1 _4980_ (.RESET_B(net277),
    .D(_0527_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .CLK(_0175_));
 sg13g2_dfrbpq_1 _4981_ (.RESET_B(net273),
    .D(_0528_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .CLK(_0176_));
 sg13g2_dfrbpq_1 _4982_ (.RESET_B(net269),
    .D(_0529_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .CLK(_0177_));
 sg13g2_dfrbpq_1 _4983_ (.RESET_B(net266),
    .D(_0530_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .CLK(_0178_));
 sg13g2_dfrbpq_1 _4984_ (.RESET_B(net262),
    .D(_0531_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .CLK(_0179_));
 sg13g2_dfrbpq_1 _4985_ (.RESET_B(net258),
    .D(_0532_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .CLK(_0180_));
 sg13g2_dfrbpq_1 _4986_ (.RESET_B(net250),
    .D(_0533_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .CLK(_0181_));
 sg13g2_dfrbpq_1 _4987_ (.RESET_B(net246),
    .D(_0534_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .CLK(_0182_));
 sg13g2_dfrbpq_1 _4988_ (.RESET_B(net242),
    .D(_0535_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .CLK(_0183_));
 sg13g2_dfrbpq_1 _4989_ (.RESET_B(net238),
    .D(_0536_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .CLK(_0184_));
 sg13g2_dfrbpq_1 _4990_ (.RESET_B(net234),
    .D(_0537_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .CLK(_0185_));
 sg13g2_dfrbpq_1 _4991_ (.RESET_B(net231),
    .D(_0538_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ),
    .CLK(_0186_));
 sg13g2_dfrbpq_1 _4992_ (.RESET_B(net227),
    .D(_0539_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .CLK(_0187_));
 sg13g2_dfrbpq_1 _4993_ (.RESET_B(net223),
    .D(_0540_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .CLK(_0188_));
 sg13g2_dfrbpq_1 _4994_ (.RESET_B(net219),
    .D(_0541_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .CLK(_0189_));
 sg13g2_dfrbpq_1 _4995_ (.RESET_B(net215),
    .D(_0542_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ),
    .CLK(_0190_));
 sg13g2_dfrbpq_1 _4996_ (.RESET_B(net211),
    .D(_0543_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .CLK(_0191_));
 sg13g2_dfrbpq_1 _4997_ (.RESET_B(net207),
    .D(_0544_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .CLK(_0192_));
 sg13g2_dfrbpq_1 _4998_ (.RESET_B(net203),
    .D(_0545_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .CLK(_0193_));
 sg13g2_dfrbpq_1 _4999_ (.RESET_B(net199),
    .D(_0546_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .CLK(_0194_));
 sg13g2_dfrbpq_1 _5000_ (.RESET_B(net195),
    .D(_0547_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .CLK(_0195_));
 sg13g2_dfrbpq_1 _5001_ (.RESET_B(net191),
    .D(_0548_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .CLK(_0196_));
 sg13g2_dfrbpq_1 _5002_ (.RESET_B(net187),
    .D(_0549_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .CLK(_0197_));
 sg13g2_dfrbpq_1 _5003_ (.RESET_B(net183),
    .D(_0550_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .CLK(_0198_));
 sg13g2_dfrbpq_1 _5004_ (.RESET_B(net179),
    .D(_0551_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .CLK(_0199_));
 sg13g2_dfrbpq_1 _5005_ (.RESET_B(net175),
    .D(_0552_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .CLK(_0200_));
 sg13g2_dfrbpq_1 _5006_ (.RESET_B(net171),
    .D(_0553_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .CLK(_0201_));
 sg13g2_dfrbpq_1 _5007_ (.RESET_B(net167),
    .D(_0554_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .CLK(_0202_));
 sg13g2_dfrbpq_1 _5008_ (.RESET_B(net163),
    .D(_0555_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ),
    .CLK(_0203_));
 sg13g2_dfrbpq_1 _5009_ (.RESET_B(net159),
    .D(_0556_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .CLK(_0204_));
 sg13g2_dfrbpq_1 _5010_ (.RESET_B(net150),
    .D(_0557_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ),
    .CLK(_0205_));
 sg13g2_dfrbpq_1 _5011_ (.RESET_B(net134),
    .D(_0558_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ),
    .CLK(_0206_));
 sg13g2_dfrbpq_1 _5012_ (.RESET_B(net126),
    .D(_0559_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .CLK(_0207_));
 sg13g2_dfrbpq_1 _5013_ (.RESET_B(net118),
    .D(_0560_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .CLK(_0208_));
 sg13g2_dfrbpq_1 _5014_ (.RESET_B(net110),
    .D(_0561_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .CLK(_0209_));
 sg13g2_dfrbpq_1 _5015_ (.RESET_B(net102),
    .D(_0562_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .CLK(_0210_));
 sg13g2_dfrbpq_1 _5016_ (.RESET_B(net94),
    .D(_0563_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .CLK(_0211_));
 sg13g2_dfrbpq_1 _5017_ (.RESET_B(net76),
    .D(_0564_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .CLK(_0212_));
 sg13g2_dfrbpq_1 _5018_ (.RESET_B(net67),
    .D(_0565_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .CLK(_0213_));
 sg13g2_dfrbpq_1 _5019_ (.RESET_B(net59),
    .D(_0566_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ),
    .CLK(_0214_));
 sg13g2_dfrbpq_1 _5020_ (.RESET_B(net51),
    .D(_0567_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .CLK(_0215_));
 sg13g2_dfrbpq_1 _5021_ (.RESET_B(net43),
    .D(_0568_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .CLK(_0216_));
 sg13g2_dfrbpq_1 _5022_ (.RESET_B(net35),
    .D(_0569_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .CLK(_0217_));
 sg13g2_dfrbpq_1 _5023_ (.RESET_B(net381),
    .D(_0570_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .CLK(_0218_));
 sg13g2_dfrbpq_1 _5024_ (.RESET_B(net373),
    .D(_0571_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .CLK(_0219_));
 sg13g2_dfrbpq_1 _5025_ (.RESET_B(net365),
    .D(_0572_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .CLK(_0220_));
 sg13g2_dfrbpq_1 _5026_ (.RESET_B(net357),
    .D(_0573_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .CLK(_0221_));
 sg13g2_dfrbpq_1 _5027_ (.RESET_B(net349),
    .D(_0574_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .CLK(_0222_));
 sg13g2_dfrbpq_1 _5028_ (.RESET_B(net318),
    .D(_0575_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .CLK(_0223_));
 sg13g2_dfrbpq_1 _5029_ (.RESET_B(net310),
    .D(_0576_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .CLK(_0224_));
 sg13g2_dfrbpq_1 _5030_ (.RESET_B(net302),
    .D(_0577_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .CLK(_0225_));
 sg13g2_dfrbpq_1 _5031_ (.RESET_B(net295),
    .D(_0578_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .CLK(_0226_));
 sg13g2_dfrbpq_1 _5032_ (.RESET_B(net287),
    .D(_0579_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .CLK(_0227_));
 sg13g2_dfrbpq_1 _5033_ (.RESET_B(net279),
    .D(_0580_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .CLK(_0228_));
 sg13g2_dfrbpq_1 _5034_ (.RESET_B(net271),
    .D(_0581_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .CLK(_0229_));
 sg13g2_dfrbpq_1 _5035_ (.RESET_B(net264),
    .D(_0582_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .CLK(_0230_));
 sg13g2_dfrbpq_1 _5036_ (.RESET_B(net252),
    .D(_0583_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .CLK(_0231_));
 sg13g2_dfrbpq_1 _5037_ (.RESET_B(net244),
    .D(_0584_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .CLK(_0232_));
 sg13g2_dfrbpq_1 _5038_ (.RESET_B(net236),
    .D(_0585_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .CLK(_0233_));
 sg13g2_dfrbpq_1 _5039_ (.RESET_B(net229),
    .D(_0586_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .CLK(_0234_));
 sg13g2_dfrbpq_1 _5040_ (.RESET_B(net221),
    .D(_0587_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .CLK(_0235_));
 sg13g2_dfrbpq_1 _5041_ (.RESET_B(net213),
    .D(_0588_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .CLK(_0236_));
 sg13g2_dfrbpq_1 _5042_ (.RESET_B(net205),
    .D(_0589_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .CLK(_0237_));
 sg13g2_dfrbpq_1 _5043_ (.RESET_B(net197),
    .D(_0590_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .CLK(_0238_));
 sg13g2_dfrbpq_1 _5044_ (.RESET_B(net189),
    .D(_0591_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .CLK(_0239_));
 sg13g2_dfrbpq_1 _5045_ (.RESET_B(net181),
    .D(_0592_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .CLK(_0240_));
 sg13g2_dfrbpq_1 _5046_ (.RESET_B(net173),
    .D(_0593_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .CLK(_0241_));
 sg13g2_dfrbpq_1 _5047_ (.RESET_B(net165),
    .D(_0594_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .CLK(_0242_));
 sg13g2_dfrbpq_1 _5048_ (.RESET_B(net157),
    .D(_0595_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .CLK(_0243_));
 sg13g2_dfrbpq_1 _5049_ (.RESET_B(net130),
    .D(_0596_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .CLK(_0244_));
 sg13g2_dfrbpq_1 _5050_ (.RESET_B(net114),
    .D(_0597_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .CLK(_0245_));
 sg13g2_dfrbpq_1 _5051_ (.RESET_B(net98),
    .D(_0598_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ),
    .CLK(_0246_));
 sg13g2_dfrbpq_1 _5052_ (.RESET_B(net72),
    .D(_0599_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .CLK(_0247_));
 sg13g2_dfrbpq_1 _5053_ (.RESET_B(net55),
    .D(_0600_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .CLK(_0248_));
 sg13g2_dfrbpq_1 _5054_ (.RESET_B(net39),
    .D(_0601_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ),
    .CLK(_0249_));
 sg13g2_dfrbpq_1 _5055_ (.RESET_B(net377),
    .D(_0602_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .CLK(_0250_));
 sg13g2_dfrbpq_1 _5056_ (.RESET_B(net361),
    .D(_0603_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .CLK(_0251_));
 sg13g2_dfrbpq_1 _5057_ (.RESET_B(net345),
    .D(_0604_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .CLK(_0252_));
 sg13g2_dfrbpq_1 _5058_ (.RESET_B(net306),
    .D(_0605_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .CLK(_0253_));
 sg13g2_dfrbpq_1 _5059_ (.RESET_B(net291),
    .D(_0606_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .CLK(_0254_));
 sg13g2_dfrbpq_1 _5060_ (.RESET_B(net275),
    .D(_0607_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ),
    .CLK(_0255_));
 sg13g2_dfrbpq_1 _5061_ (.RESET_B(net260),
    .D(_0608_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .CLK(_0256_));
 sg13g2_dfrbpq_1 _5062_ (.RESET_B(net240),
    .D(_0609_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .CLK(_0257_));
 sg13g2_dfrbpq_1 _5063_ (.RESET_B(net225),
    .D(_0610_),
    .Q(\blue_tmds_par[0] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _5064_ (.RESET_B(net217),
    .D(_0611_),
    .Q(\blue_tmds_par[1] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _5065_ (.RESET_B(net209),
    .D(_0612_),
    .Q(\blue_tmds_par[2] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _5066_ (.RESET_B(net201),
    .D(_0613_),
    .Q(\blue_tmds_par[3] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _5067_ (.RESET_B(net193),
    .D(_0614_),
    .Q(\blue_tmds_par[5] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _5068_ (.RESET_B(net185),
    .D(_0615_),
    .Q(\blue_tmds_par[6] ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _5069_ (.RESET_B(net177),
    .D(_0616_),
    .Q(\blue_tmds_par[7] ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _5070_ (.RESET_B(net169),
    .D(_0617_),
    .Q(\blue_tmds_par[8] ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _5071_ (.RESET_B(net161),
    .D(_0618_),
    .Q(\blue_tmds_par[9] ),
    .CLK(net641));
 sg13g2_dfrbpq_2 _5072_ (.RESET_B(net146),
    .D(_0619_),
    .Q(\tmds_green.dc_balancing_reg[1] ),
    .CLK(net648));
 sg13g2_dfrbpq_1 _5073_ (.RESET_B(net122),
    .D(_0620_),
    .Q(\tmds_green.dc_balancing_reg[2] ),
    .CLK(net648));
 sg13g2_dfrbpq_1 _5074_ (.RESET_B(net106),
    .D(_0621_),
    .Q(\tmds_green.dc_balancing_reg[3] ),
    .CLK(net648));
 sg13g2_dfrbpq_2 _5075_ (.RESET_B(net90),
    .D(_0622_),
    .Q(\tmds_green.dc_balancing_reg[4] ),
    .CLK(net648));
 sg13g2_dfrbpq_1 _5076_ (.RESET_B(net63),
    .D(net407),
    .Q(\clockdiv.q0 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _5077_ (.RESET_B(net47),
    .D(_0624_),
    .Q(\tmds_blue.dc_balancing_reg[1] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _5078_ (.RESET_B(net31),
    .D(_0625_),
    .Q(\tmds_blue.dc_balancing_reg[2] ),
    .CLK(net641));
 sg13g2_dfrbpq_2 _5079_ (.RESET_B(net369),
    .D(_0626_),
    .Q(\tmds_blue.dc_balancing_reg[3] ),
    .CLK(net643));
 sg13g2_dfrbpq_2 _5080_ (.RESET_B(net353),
    .D(_0627_),
    .Q(\tmds_blue.dc_balancing_reg[4] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _5081_ (.RESET_B(net314),
    .D(_0628_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .CLK(_0258_));
 sg13g2_dfrbpq_1 _5082_ (.RESET_B(net283),
    .D(_0629_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .CLK(_0259_));
 sg13g2_dfrbpq_1 _5083_ (.RESET_B(net248),
    .D(_0630_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .CLK(_0260_));
 sg13g2_dfrbpq_1 _5084_ (.RESET_B(net403),
    .D(_0631_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .CLK(_0261_));
 sg13g2_dfrbpq_1 _5085_ (.RESET_B(net799),
    .D(\serialize.n428[0] ),
    .Q(\serialize.n453 ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5086_ (.RESET_B(net799),
    .D(\serialize.n428[1] ),
    .Q(\serialize.n455 ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5087_ (.RESET_B(net799),
    .D(\serialize.n428[2] ),
    .Q(\serialize.n414[0] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5088_ (.RESET_B(net801),
    .D(\serialize.n428[3] ),
    .Q(\serialize.n414[1] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5089_ (.RESET_B(net798),
    .D(\serialize.n428[4] ),
    .Q(\serialize.n414[2] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5090_ (.RESET_B(net801),
    .D(\serialize.n428[5] ),
    .Q(\serialize.n414[3] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5091_ (.RESET_B(net798),
    .D(net428),
    .Q(\serialize.n414[4] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5092_ (.RESET_B(net801),
    .D(\serialize.n428[7] ),
    .Q(\serialize.n414[5] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5093_ (.RESET_B(net798),
    .D(\serialize.n428[8] ),
    .Q(\serialize.n414[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5094_ (.RESET_B(net801),
    .D(\serialize.n428[9] ),
    .Q(\serialize.n414[7] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5095_ (.RESET_B(net801),
    .D(\serialize.n431[0] ),
    .Q(\serialize.n459 ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5096_ (.RESET_B(net801),
    .D(\serialize.n431[1] ),
    .Q(\serialize.n461 ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5097_ (.RESET_B(net801),
    .D(\serialize.n431[2] ),
    .Q(\serialize.n420[0] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5098_ (.RESET_B(net801),
    .D(\serialize.n431[3] ),
    .Q(\serialize.n420[1] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5099_ (.RESET_B(net800),
    .D(\serialize.n431[4] ),
    .Q(\serialize.n420[2] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5100_ (.RESET_B(net800),
    .D(\serialize.n431[5] ),
    .Q(\serialize.n420[3] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5101_ (.RESET_B(net800),
    .D(net416),
    .Q(\serialize.n420[4] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5102_ (.RESET_B(net797),
    .D(net695),
    .Q(\serialize.n420[6] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5103_ (.RESET_B(net800),
    .D(\serialize.n429[0] ),
    .Q(\serialize.n456 ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5104_ (.RESET_B(net800),
    .D(\serialize.n429[1] ),
    .Q(\serialize.n458 ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5105_ (.RESET_B(net800),
    .D(\serialize.n429[2] ),
    .Q(\serialize.n417[0] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5106_ (.RESET_B(net800),
    .D(\serialize.n429[3] ),
    .Q(\serialize.n417[1] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5107_ (.RESET_B(net796),
    .D(\serialize.n429[4] ),
    .Q(\serialize.n417[2] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5108_ (.RESET_B(net800),
    .D(\serialize.n429[5] ),
    .Q(\serialize.n417[3] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5109_ (.RESET_B(net796),
    .D(\serialize.n429[6] ),
    .Q(\serialize.n417[4] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5110_ (.RESET_B(net796),
    .D(\serialize.n429[7] ),
    .Q(\serialize.n417[5] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5111_ (.RESET_B(net796),
    .D(\serialize.n429[8] ),
    .Q(\serialize.n417[6] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5112_ (.RESET_B(net797),
    .D(\serialize.n429[9] ),
    .Q(\serialize.n417[7] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _5113_ (.RESET_B(net796),
    .D(\serialize.n433[0] ),
    .Q(\serialize.bit_cnt[0] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _5114_ (.RESET_B(net796),
    .D(\serialize.n433[1] ),
    .Q(\serialize.bit_cnt[1] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5115_ (.RESET_B(net796),
    .D(_0262_),
    .Q(_0004_),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5116_ (.RESET_B(net799),
    .D(\serialize.n427[0] ),
    .Q(\serialize.n450 ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5117_ (.RESET_B(net799),
    .D(\serialize.n427[1] ),
    .Q(\serialize.n452 ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5118_ (.RESET_B(net799),
    .D(\serialize.n427[2] ),
    .Q(\serialize.n411[0] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5119_ (.RESET_B(net799),
    .D(\serialize.n427[3] ),
    .Q(\serialize.n411[1] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5120_ (.RESET_B(net798),
    .D(\serialize.n427[4] ),
    .Q(\serialize.n411[2] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5121_ (.RESET_B(net799),
    .D(\serialize.n427[5] ),
    .Q(\serialize.n411[3] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5122_ (.RESET_B(net798),
    .D(net420),
    .Q(\serialize.n411[4] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5123_ (.RESET_B(net798),
    .D(\serialize.n427[7] ),
    .Q(\serialize.n411[5] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5124_ (.RESET_B(net798),
    .D(\serialize.n427[8] ),
    .Q(\serialize.n411[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5125_ (.RESET_B(net798),
    .D(\serialize.n427[9] ),
    .Q(\serialize.n411[7] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_tiehi _4785__32 (.L_HI(net32));
 sg13g2_tiehi _4949__33 (.L_HI(net33));
 sg13g2_tiehi _4784__34 (.L_HI(net34));
 sg13g2_tiehi _5022__35 (.L_HI(net35));
 sg13g2_tiehi _4783__36 (.L_HI(net36));
 sg13g2_tiehi _4948__37 (.L_HI(net37));
 sg13g2_tiehi _4782__38 (.L_HI(net38));
 sg13g2_tiehi _5054__39 (.L_HI(net39));
 sg13g2_tiehi _4781__40 (.L_HI(net40));
 sg13g2_tiehi _4947__41 (.L_HI(net41));
 sg13g2_tiehi _4780__42 (.L_HI(net42));
 sg13g2_tiehi _5021__43 (.L_HI(net43));
 sg13g2_tiehi _4779__44 (.L_HI(net44));
 sg13g2_tiehi _4946__45 (.L_HI(net45));
 sg13g2_tiehi _4778__46 (.L_HI(net46));
 sg13g2_tiehi _5077__47 (.L_HI(net47));
 sg13g2_tiehi _4777__48 (.L_HI(net48));
 sg13g2_tiehi _4945__49 (.L_HI(net49));
 sg13g2_tiehi _4776__50 (.L_HI(net50));
 sg13g2_tiehi _5020__51 (.L_HI(net51));
 sg13g2_tiehi _4775__52 (.L_HI(net52));
 sg13g2_tiehi _4944__53 (.L_HI(net53));
 sg13g2_tiehi _4774__54 (.L_HI(net54));
 sg13g2_tiehi _5053__55 (.L_HI(net55));
 sg13g2_tiehi _4773__56 (.L_HI(net56));
 sg13g2_tiehi _4943__57 (.L_HI(net57));
 sg13g2_tiehi _4772__58 (.L_HI(net58));
 sg13g2_tiehi _5019__59 (.L_HI(net59));
 sg13g2_tiehi _4771__60 (.L_HI(net60));
 sg13g2_tiehi _4942__61 (.L_HI(net61));
 sg13g2_tiehi _4770__62 (.L_HI(net62));
 sg13g2_tiehi _5076__63 (.L_HI(net63));
 sg13g2_tiehi _4769__64 (.L_HI(net64));
 sg13g2_tiehi _4941__65 (.L_HI(net65));
 sg13g2_tiehi _4768__66 (.L_HI(net66));
 sg13g2_tiehi _5018__67 (.L_HI(net67));
 sg13g2_tiehi _4767__68 (.L_HI(net68));
 sg13g2_tiehi _4766__69 (.L_HI(net69));
 sg13g2_tiehi _4940__70 (.L_HI(net70));
 sg13g2_tiehi _4765__71 (.L_HI(net71));
 sg13g2_tiehi _5052__72 (.L_HI(net72));
 sg13g2_tiehi _4764__73 (.L_HI(net73));
 sg13g2_tiehi _4939__74 (.L_HI(net74));
 sg13g2_tiehi _4763__75 (.L_HI(net75));
 sg13g2_tiehi _5017__76 (.L_HI(net76));
 sg13g2_tiehi _4762__77 (.L_HI(net77));
 sg13g2_tiehi _4761__78 (.L_HI(net78));
 sg13g2_tiehi _4760__79 (.L_HI(net79));
 sg13g2_tiehi _4759__80 (.L_HI(net80));
 sg13g2_tiehi _4758__81 (.L_HI(net81));
 sg13g2_tiehi _4757__82 (.L_HI(net82));
 sg13g2_tiehi _4756__83 (.L_HI(net83));
 sg13g2_tiehi _4755__84 (.L_HI(net84));
 sg13g2_tiehi _4754__85 (.L_HI(net85));
 sg13g2_tiehi _4753__86 (.L_HI(net86));
 sg13g2_tiehi _4752__87 (.L_HI(net87));
 sg13g2_tiehi _4938__88 (.L_HI(net88));
 sg13g2_tiehi _4751__89 (.L_HI(net89));
 sg13g2_tiehi _5075__90 (.L_HI(net90));
 sg13g2_tiehi _4750__91 (.L_HI(net91));
 sg13g2_tiehi _4937__92 (.L_HI(net92));
 sg13g2_tiehi _4749__93 (.L_HI(net93));
 sg13g2_tiehi _5016__94 (.L_HI(net94));
 sg13g2_tiehi _4748__95 (.L_HI(net95));
 sg13g2_tiehi _4932__96 (.L_HI(net96));
 sg13g2_tiehi _4747__97 (.L_HI(net97));
 sg13g2_tiehi _5051__98 (.L_HI(net98));
 sg13g2_tiehi _4746__99 (.L_HI(net99));
 sg13g2_tiehi _4931__100 (.L_HI(net100));
 sg13g2_tiehi _4745__101 (.L_HI(net101));
 sg13g2_tiehi _5015__102 (.L_HI(net102));
 sg13g2_tiehi _4744__103 (.L_HI(net103));
 sg13g2_tiehi _4930__104 (.L_HI(net104));
 sg13g2_tiehi _4743__105 (.L_HI(net105));
 sg13g2_tiehi _5074__106 (.L_HI(net106));
 sg13g2_tiehi _4742__107 (.L_HI(net107));
 sg13g2_tiehi _4929__108 (.L_HI(net108));
 sg13g2_tiehi _4741__109 (.L_HI(net109));
 sg13g2_tiehi _5014__110 (.L_HI(net110));
 sg13g2_tiehi _4740__111 (.L_HI(net111));
 sg13g2_tiehi _4928__112 (.L_HI(net112));
 sg13g2_tiehi _4739__113 (.L_HI(net113));
 sg13g2_tiehi _5050__114 (.L_HI(net114));
 sg13g2_tiehi _4738__115 (.L_HI(net115));
 sg13g2_tiehi _4927__116 (.L_HI(net116));
 sg13g2_tiehi _4737__117 (.L_HI(net117));
 sg13g2_tiehi _5013__118 (.L_HI(net118));
 sg13g2_tiehi _4736__119 (.L_HI(net119));
 sg13g2_tiehi _4926__120 (.L_HI(net120));
 sg13g2_tiehi _4735__121 (.L_HI(net121));
 sg13g2_tiehi _5073__122 (.L_HI(net122));
 sg13g2_tiehi _4734__123 (.L_HI(net123));
 sg13g2_tiehi _4925__124 (.L_HI(net124));
 sg13g2_tiehi _4733__125 (.L_HI(net125));
 sg13g2_tiehi _5012__126 (.L_HI(net126));
 sg13g2_tiehi _4732__127 (.L_HI(net127));
 sg13g2_tiehi _4924__128 (.L_HI(net128));
 sg13g2_tiehi _4731__129 (.L_HI(net129));
 sg13g2_tiehi _5049__130 (.L_HI(net130));
 sg13g2_tiehi _4730__131 (.L_HI(net131));
 sg13g2_tiehi _4923__132 (.L_HI(net132));
 sg13g2_tiehi _4729__133 (.L_HI(net133));
 sg13g2_tiehi _5011__134 (.L_HI(net134));
 sg13g2_tiehi _4728__135 (.L_HI(net135));
 sg13g2_tiehi _4727__136 (.L_HI(net136));
 sg13g2_tiehi _4726__137 (.L_HI(net137));
 sg13g2_tiehi _4725__138 (.L_HI(net138));
 sg13g2_tiehi _4724__139 (.L_HI(net139));
 sg13g2_tiehi _4723__140 (.L_HI(net140));
 sg13g2_tiehi _4722__141 (.L_HI(net141));
 sg13g2_tiehi _4721__142 (.L_HI(net142));
 sg13g2_tiehi _4720__143 (.L_HI(net143));
 sg13g2_tiehi _4922__144 (.L_HI(net144));
 sg13g2_tiehi _4719__145 (.L_HI(net145));
 sg13g2_tiehi _5072__146 (.L_HI(net146));
 sg13g2_tiehi _4718__147 (.L_HI(net147));
 sg13g2_tiehi _4921__148 (.L_HI(net148));
 sg13g2_tiehi _4717__149 (.L_HI(net149));
 sg13g2_tiehi _5010__150 (.L_HI(net150));
 sg13g2_tiehi _4716__151 (.L_HI(net151));
 sg13g2_tiehi _4715__152 (.L_HI(net152));
 sg13g2_tiehi _4714__153 (.L_HI(net153));
 sg13g2_tiehi _4713__154 (.L_HI(net154));
 sg13g2_tiehi _4920__155 (.L_HI(net155));
 sg13g2_tiehi _4712__156 (.L_HI(net156));
 sg13g2_tiehi _5048__157 (.L_HI(net157));
 sg13g2_tiehi _4919__158 (.L_HI(net158));
 sg13g2_tiehi _5009__159 (.L_HI(net159));
 sg13g2_tiehi _4918__160 (.L_HI(net160));
 sg13g2_tiehi _5071__161 (.L_HI(net161));
 sg13g2_tiehi _4917__162 (.L_HI(net162));
 sg13g2_tiehi _5008__163 (.L_HI(net163));
 sg13g2_tiehi _4916__164 (.L_HI(net164));
 sg13g2_tiehi _5047__165 (.L_HI(net165));
 sg13g2_tiehi _4915__166 (.L_HI(net166));
 sg13g2_tiehi _5007__167 (.L_HI(net167));
 sg13g2_tiehi _4914__168 (.L_HI(net168));
 sg13g2_tiehi _5070__169 (.L_HI(net169));
 sg13g2_tiehi _4913__170 (.L_HI(net170));
 sg13g2_tiehi _5006__171 (.L_HI(net171));
 sg13g2_tiehi _4912__172 (.L_HI(net172));
 sg13g2_tiehi _5046__173 (.L_HI(net173));
 sg13g2_tiehi _4911__174 (.L_HI(net174));
 sg13g2_tiehi _5005__175 (.L_HI(net175));
 sg13g2_tiehi _4910__176 (.L_HI(net176));
 sg13g2_tiehi _5069__177 (.L_HI(net177));
 sg13g2_tiehi _4909__178 (.L_HI(net178));
 sg13g2_tiehi _5004__179 (.L_HI(net179));
 sg13g2_tiehi _4908__180 (.L_HI(net180));
 sg13g2_tiehi _5045__181 (.L_HI(net181));
 sg13g2_tiehi _4907__182 (.L_HI(net182));
 sg13g2_tiehi _5003__183 (.L_HI(net183));
 sg13g2_tiehi _4906__184 (.L_HI(net184));
 sg13g2_tiehi _5068__185 (.L_HI(net185));
 sg13g2_tiehi _4905__186 (.L_HI(net186));
 sg13g2_tiehi _5002__187 (.L_HI(net187));
 sg13g2_tiehi _4904__188 (.L_HI(net188));
 sg13g2_tiehi _5044__189 (.L_HI(net189));
 sg13g2_tiehi _4903__190 (.L_HI(net190));
 sg13g2_tiehi _5001__191 (.L_HI(net191));
 sg13g2_tiehi _4902__192 (.L_HI(net192));
 sg13g2_tiehi _5067__193 (.L_HI(net193));
 sg13g2_tiehi _4901__194 (.L_HI(net194));
 sg13g2_tiehi _5000__195 (.L_HI(net195));
 sg13g2_tiehi _4900__196 (.L_HI(net196));
 sg13g2_tiehi _5043__197 (.L_HI(net197));
 sg13g2_tiehi _4899__198 (.L_HI(net198));
 sg13g2_tiehi _4999__199 (.L_HI(net199));
 sg13g2_tiehi _4898__200 (.L_HI(net200));
 sg13g2_tiehi _5066__201 (.L_HI(net201));
 sg13g2_tiehi _4897__202 (.L_HI(net202));
 sg13g2_tiehi _4998__203 (.L_HI(net203));
 sg13g2_tiehi _4896__204 (.L_HI(net204));
 sg13g2_tiehi _5042__205 (.L_HI(net205));
 sg13g2_tiehi _4895__206 (.L_HI(net206));
 sg13g2_tiehi _4997__207 (.L_HI(net207));
 sg13g2_tiehi _4894__208 (.L_HI(net208));
 sg13g2_tiehi _5065__209 (.L_HI(net209));
 sg13g2_tiehi _4893__210 (.L_HI(net210));
 sg13g2_tiehi _4996__211 (.L_HI(net211));
 sg13g2_tiehi _4892__212 (.L_HI(net212));
 sg13g2_tiehi _5041__213 (.L_HI(net213));
 sg13g2_tiehi _4891__214 (.L_HI(net214));
 sg13g2_tiehi _4995__215 (.L_HI(net215));
 sg13g2_tiehi _4890__216 (.L_HI(net216));
 sg13g2_tiehi _5064__217 (.L_HI(net217));
 sg13g2_tiehi _4889__218 (.L_HI(net218));
 sg13g2_tiehi _4994__219 (.L_HI(net219));
 sg13g2_tiehi _4888__220 (.L_HI(net220));
 sg13g2_tiehi _5040__221 (.L_HI(net221));
 sg13g2_tiehi _4887__222 (.L_HI(net222));
 sg13g2_tiehi _4993__223 (.L_HI(net223));
 sg13g2_tiehi _4886__224 (.L_HI(net224));
 sg13g2_tiehi _5063__225 (.L_HI(net225));
 sg13g2_tiehi _4885__226 (.L_HI(net226));
 sg13g2_tiehi _4992__227 (.L_HI(net227));
 sg13g2_tiehi _4884__228 (.L_HI(net228));
 sg13g2_tiehi _5039__229 (.L_HI(net229));
 sg13g2_tiehi _4883__230 (.L_HI(net230));
 sg13g2_tiehi _4991__231 (.L_HI(net231));
 sg13g2_tiehi _4882__232 (.L_HI(net232));
 sg13g2_tiehi _4881__233 (.L_HI(net233));
 sg13g2_tiehi _4990__234 (.L_HI(net234));
 sg13g2_tiehi _4880__235 (.L_HI(net235));
 sg13g2_tiehi _5038__236 (.L_HI(net236));
 sg13g2_tiehi _4879__237 (.L_HI(net237));
 sg13g2_tiehi _4989__238 (.L_HI(net238));
 sg13g2_tiehi _4878__239 (.L_HI(net239));
 sg13g2_tiehi _5062__240 (.L_HI(net240));
 sg13g2_tiehi _4877__241 (.L_HI(net241));
 sg13g2_tiehi _4988__242 (.L_HI(net242));
 sg13g2_tiehi _4876__243 (.L_HI(net243));
 sg13g2_tiehi _5037__244 (.L_HI(net244));
 sg13g2_tiehi _4875__245 (.L_HI(net245));
 sg13g2_tiehi _4987__246 (.L_HI(net246));
 sg13g2_tiehi _4874__247 (.L_HI(net247));
 sg13g2_tiehi _5083__248 (.L_HI(net248));
 sg13g2_tiehi _4873__249 (.L_HI(net249));
 sg13g2_tiehi _4986__250 (.L_HI(net250));
 sg13g2_tiehi _4872__251 (.L_HI(net251));
 sg13g2_tiehi _5036__252 (.L_HI(net252));
 sg13g2_tiehi _4711__253 (.L_HI(net253));
 sg13g2_tiehi _4933__254 (.L_HI(net254));
 sg13g2_tiehi _4934__255 (.L_HI(net255));
 sg13g2_tiehi _4935__256 (.L_HI(net256));
 sg13g2_tiehi _4871__257 (.L_HI(net257));
 sg13g2_tiehi _4985__258 (.L_HI(net258));
 sg13g2_tiehi _4870__259 (.L_HI(net259));
 sg13g2_tiehi _5061__260 (.L_HI(net260));
 sg13g2_tiehi _4869__261 (.L_HI(net261));
 sg13g2_tiehi _4984__262 (.L_HI(net262));
 sg13g2_tiehi _4868__263 (.L_HI(net263));
 sg13g2_tiehi _5035__264 (.L_HI(net264));
 sg13g2_tiehi _4867__265 (.L_HI(net265));
 sg13g2_tiehi _4983__266 (.L_HI(net266));
 sg13g2_tiehi _4866__267 (.L_HI(net267));
 sg13g2_tiehi _4865__268 (.L_HI(net268));
 sg13g2_tiehi _4982__269 (.L_HI(net269));
 sg13g2_tiehi _4864__270 (.L_HI(net270));
 sg13g2_tiehi _5034__271 (.L_HI(net271));
 sg13g2_tiehi _4863__272 (.L_HI(net272));
 sg13g2_tiehi _4981__273 (.L_HI(net273));
 sg13g2_tiehi _4862__274 (.L_HI(net274));
 sg13g2_tiehi _5060__275 (.L_HI(net275));
 sg13g2_tiehi _4861__276 (.L_HI(net276));
 sg13g2_tiehi _4980__277 (.L_HI(net277));
 sg13g2_tiehi _4860__278 (.L_HI(net278));
 sg13g2_tiehi _5033__279 (.L_HI(net279));
 sg13g2_tiehi _4859__280 (.L_HI(net280));
 sg13g2_tiehi _4979__281 (.L_HI(net281));
 sg13g2_tiehi _4858__282 (.L_HI(net282));
 sg13g2_tiehi _5082__283 (.L_HI(net283));
 sg13g2_tiehi _4857__284 (.L_HI(net284));
 sg13g2_tiehi _4978__285 (.L_HI(net285));
 sg13g2_tiehi _4856__286 (.L_HI(net286));
 sg13g2_tiehi _5032__287 (.L_HI(net287));
 sg13g2_tiehi _4855__288 (.L_HI(net288));
 sg13g2_tiehi _4977__289 (.L_HI(net289));
 sg13g2_tiehi _4854__290 (.L_HI(net290));
 sg13g2_tiehi _5059__291 (.L_HI(net291));
 sg13g2_tiehi _4853__292 (.L_HI(net292));
 sg13g2_tiehi _4976__293 (.L_HI(net293));
 sg13g2_tiehi _4852__294 (.L_HI(net294));
 sg13g2_tiehi _5031__295 (.L_HI(net295));
 sg13g2_tiehi _4851__296 (.L_HI(net296));
 sg13g2_tiehi _4975__297 (.L_HI(net297));
 sg13g2_tiehi _4850__298 (.L_HI(net298));
 sg13g2_tiehi _4849__299 (.L_HI(net299));
 sg13g2_tiehi _4974__300 (.L_HI(net300));
 sg13g2_tiehi _4848__301 (.L_HI(net301));
 sg13g2_tiehi _5030__302 (.L_HI(net302));
 sg13g2_tiehi _4847__303 (.L_HI(net303));
 sg13g2_tiehi _4973__304 (.L_HI(net304));
 sg13g2_tiehi _4846__305 (.L_HI(net305));
 sg13g2_tiehi _5058__306 (.L_HI(net306));
 sg13g2_tiehi _4845__307 (.L_HI(net307));
 sg13g2_tiehi _4972__308 (.L_HI(net308));
 sg13g2_tiehi _4844__309 (.L_HI(net309));
 sg13g2_tiehi _5029__310 (.L_HI(net310));
 sg13g2_tiehi _4843__311 (.L_HI(net311));
 sg13g2_tiehi _4971__312 (.L_HI(net312));
 sg13g2_tiehi _4842__313 (.L_HI(net313));
 sg13g2_tiehi _5081__314 (.L_HI(net314));
 sg13g2_tiehi _4841__315 (.L_HI(net315));
 sg13g2_tiehi _4970__316 (.L_HI(net316));
 sg13g2_tiehi _4840__317 (.L_HI(net317));
 sg13g2_tiehi _5028__318 (.L_HI(net318));
 sg13g2_tiehi _4839__319 (.L_HI(net319));
 sg13g2_tiehi _4969__320 (.L_HI(net320));
 sg13g2_tiehi _4838__321 (.L_HI(net321));
 sg13g2_tiehi _4837__322 (.L_HI(net322));
 sg13g2_tiehi _4836__323 (.L_HI(net323));
 sg13g2_tiehi _4835__324 (.L_HI(net324));
 sg13g2_tiehi _4834__325 (.L_HI(net325));
 sg13g2_tiehi _4833__326 (.L_HI(net326));
 sg13g2_tiehi _4832__327 (.L_HI(net327));
 sg13g2_tiehi _4831__328 (.L_HI(net328));
 sg13g2_tiehi _4830__329 (.L_HI(net329));
 sg13g2_tiehi _4829__330 (.L_HI(net330));
 sg13g2_tiehi _4828__331 (.L_HI(net331));
 sg13g2_tiehi _4827__332 (.L_HI(net332));
 sg13g2_tiehi _4826__333 (.L_HI(net333));
 sg13g2_tiehi _4825__334 (.L_HI(net334));
 sg13g2_tiehi _4824__335 (.L_HI(net335));
 sg13g2_tiehi _4823__336 (.L_HI(net336));
 sg13g2_tiehi _4822__337 (.L_HI(net337));
 sg13g2_tiehi _4821__338 (.L_HI(net338));
 sg13g2_tiehi _4820__339 (.L_HI(net339));
 sg13g2_tiehi _4819__340 (.L_HI(net340));
 sg13g2_tiehi _4818__341 (.L_HI(net341));
 sg13g2_tiehi _4817__342 (.L_HI(net342));
 sg13g2_tiehi _4816__343 (.L_HI(net343));
 sg13g2_tiehi _4815__344 (.L_HI(net344));
 sg13g2_tiehi _5057__345 (.L_HI(net345));
 sg13g2_tiehi _4814__346 (.L_HI(net346));
 sg13g2_tiehi _4968__347 (.L_HI(net347));
 sg13g2_tiehi _4813__348 (.L_HI(net348));
 sg13g2_tiehi _5027__349 (.L_HI(net349));
 sg13g2_tiehi _4812__350 (.L_HI(net350));
 sg13g2_tiehi _4967__351 (.L_HI(net351));
 sg13g2_tiehi _4811__352 (.L_HI(net352));
 sg13g2_tiehi _5080__353 (.L_HI(net353));
 sg13g2_tiehi _4810__354 (.L_HI(net354));
 sg13g2_tiehi _4966__355 (.L_HI(net355));
 sg13g2_tiehi _4809__356 (.L_HI(net356));
 sg13g2_tiehi _5026__357 (.L_HI(net357));
 sg13g2_tiehi _4808__358 (.L_HI(net358));
 sg13g2_tiehi _4965__359 (.L_HI(net359));
 sg13g2_tiehi _4807__360 (.L_HI(net360));
 sg13g2_tiehi _5056__361 (.L_HI(net361));
 sg13g2_tiehi _4806__362 (.L_HI(net362));
 sg13g2_tiehi _4964__363 (.L_HI(net363));
 sg13g2_tiehi _4805__364 (.L_HI(net364));
 sg13g2_tiehi _5025__365 (.L_HI(net365));
 sg13g2_tiehi _4804__366 (.L_HI(net366));
 sg13g2_tiehi _4963__367 (.L_HI(net367));
 sg13g2_tiehi _4803__368 (.L_HI(net368));
 sg13g2_tiehi _5079__369 (.L_HI(net369));
 sg13g2_tiehi _4802__370 (.L_HI(net370));
 sg13g2_tiehi _4962__371 (.L_HI(net371));
 sg13g2_tiehi _4801__372 (.L_HI(net372));
 sg13g2_tiehi _5024__373 (.L_HI(net373));
 sg13g2_tiehi _4800__374 (.L_HI(net374));
 sg13g2_tiehi _4961__375 (.L_HI(net375));
 sg13g2_tiehi _4799__376 (.L_HI(net376));
 sg13g2_tiehi _5055__377 (.L_HI(net377));
 sg13g2_tiehi _4798__378 (.L_HI(net378));
 sg13g2_tiehi _4960__379 (.L_HI(net379));
 sg13g2_tiehi _4797__380 (.L_HI(net380));
 sg13g2_tiehi _5023__381 (.L_HI(net381));
 sg13g2_tiehi _4796__382 (.L_HI(net382));
 sg13g2_tiehi _4959__383 (.L_HI(net383));
 sg13g2_tiehi _4795__384 (.L_HI(net384));
 sg13g2_tiehi _4958__385 (.L_HI(net385));
 sg13g2_tiehi _4794__386 (.L_HI(net386));
 sg13g2_tiehi _4957__387 (.L_HI(net387));
 sg13g2_tiehi _4793__388 (.L_HI(net388));
 sg13g2_tiehi _4956__389 (.L_HI(net389));
 sg13g2_tiehi _4792__390 (.L_HI(net390));
 sg13g2_tiehi _4955__391 (.L_HI(net391));
 sg13g2_tiehi _4791__392 (.L_HI(net392));
 sg13g2_tiehi _4954__393 (.L_HI(net393));
 sg13g2_tiehi _4790__394 (.L_HI(net394));
 sg13g2_tiehi _4953__395 (.L_HI(net395));
 sg13g2_tiehi _4789__396 (.L_HI(net396));
 sg13g2_tiehi _4952__397 (.L_HI(net397));
 sg13g2_tiehi _4788__398 (.L_HI(net398));
 sg13g2_tiehi _4951__399 (.L_HI(net399));
 sg13g2_tiehi _4787__400 (.L_HI(net400));
 sg13g2_tiehi _4950__401 (.L_HI(net401));
 sg13g2_tiehi _4936__402 (.L_HI(net402));
 sg13g2_tiehi _5084__403 (.L_HI(net403));
 sg13g2_tiehi _4786__404 (.L_HI(net404));
 sg13g2_inv_1 _2537__1 (.Y(net405),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo heichips25_bagel_22 (.L_LO(net22));
 sg13g2_tielo heichips25_bagel_23 (.L_LO(net23));
 sg13g2_tielo heichips25_bagel_24 (.L_LO(net24));
 sg13g2_tielo heichips25_bagel_25 (.L_LO(net25));
 sg13g2_tielo heichips25_bagel_26 (.L_LO(net26));
 sg13g2_tielo heichips25_bagel_27 (.L_LO(net27));
 sg13g2_tielo heichips25_bagel_28 (.L_LO(net28));
 sg13g2_tielo heichips25_bagel_29 (.L_LO(net29));
 sg13g2_tielo heichips25_bagel_30 (.L_LO(net30));
 sg13g2_tiehi _5078__31 (.L_HI(net31));
 sg13g2_buf_8 _5510_ (.A(\videogen.mem_row ),
    .X(net11));
 sg13g2_buf_1 _5511_ (.A(net600),
    .X(net12));
 sg13g2_buf_8 fanout542 (.A(_1111_),
    .X(net542));
 sg13g2_buf_8 fanout543 (.A(_0673_),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(_1055_),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(_1021_),
    .X(net545));
 sg13g2_buf_8 fanout546 (.A(_1031_),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(_1176_),
    .X(net547));
 sg13g2_buf_8 fanout548 (.A(_0855_),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(net558),
    .X(net549));
 sg13g2_buf_1 fanout550 (.A(net558),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(net558),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net557),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net557),
    .X(net554));
 sg13g2_buf_8 fanout555 (.A(net557),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(_1255_),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(net568),
    .X(net559));
 sg13g2_buf_1 fanout560 (.A(net568),
    .X(net560));
 sg13g2_buf_8 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_8 fanout562 (.A(net568),
    .X(net562));
 sg13g2_buf_8 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(net567),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_8 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(_1253_),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(net571),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_8 fanout571 (.A(_0837_),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(net576),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(net576),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(_0690_),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(net581),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net581),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(_0690_),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(net591),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net591),
    .X(net584));
 sg13g2_buf_8 fanout585 (.A(net591),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(net590),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(net590),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(_0675_),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(net595),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(_0639_),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(net599),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(net599),
    .X(net597));
 sg13g2_buf_1 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(_0638_),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(\videogen.mem_read ),
    .X(net600));
 sg13g2_buf_8 fanout601 (.A(\tmds_green.n132 ),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(\tmds_green.n100 ),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(\tmds_blue.n100 ),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(display_enable),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(\videogen.fancy_shader.video_y[1] ),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(\videogen.fancy_shader.video_y[0] ),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(\videogen.fancy_shader.n646[8] ),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(\videogen.fancy_shader.n646[3] ),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_8 fanout613 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(net623),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net623),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(net628),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(\videogen.fancy_shader.video_x[7] ),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(\videogen.fancy_shader.video_x[0] ),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net650),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net639),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net639),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net639),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net650),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net650),
    .X(net643));
 sg13g2_buf_8 fanout644 (.A(net646),
    .X(net644));
 sg13g2_buf_1 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net649),
    .X(net646));
 sg13g2_buf_8 fanout647 (.A(net649),
    .X(net647));
 sg13g2_buf_1 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(clk_video),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net656),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(net655),
    .X(net653));
 sg13g2_buf_1 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net694),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(net660),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(net660),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(net694),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(net663),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net673),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(net667),
    .X(net664));
 sg13g2_buf_1 fanout665 (.A(net667),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net673),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net673),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net673),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net672),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_8 fanout673 (.A(net694),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net678),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(net678),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net678),
    .X(net676));
 sg13g2_buf_1 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_8 fanout678 (.A(net683),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(net683),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(net694),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net693),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(net693),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net693),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(net692),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(\clockdiv.q2temp ),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net430),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(net701),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net701),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net701),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(\serialize.n410 ),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(net707),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net706),
    .X(net704));
 sg13g2_buf_1 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net746),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(net711),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(net711),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(net746),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(net714),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(net724),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(net718),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(net718),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(net724),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(net724),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net746),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net734),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(net734),
    .X(net728));
 sg13g2_buf_1 fanout729 (.A(net734),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net734),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net746),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(net739),
    .X(net735));
 sg13g2_buf_1 fanout736 (.A(net739),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net745),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net745),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(net745),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(net745),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(\clockdiv.q1 ),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(net749),
    .X(net747));
 sg13g2_buf_1 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(_0648_),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(_0648_),
    .X(net751));
 sg13g2_buf_8 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net761),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(net761),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(net760),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net760),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(ui_in[7]),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net766),
    .X(net762));
 sg13g2_buf_1 fanout763 (.A(net766),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(ui_in[6]),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net771),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_8 fanout771 (.A(ui_in[6]),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net776),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_8 fanout776 (.A(ui_in[5]),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net781),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(net781),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net781),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(ui_in[5]),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net792),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net792),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net786),
    .X(net784));
 sg13g2_buf_1 fanout785 (.A(net786),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net792),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net791),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net791),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net791),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(ui_in[4]),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(rst_n),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net803),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net803),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(net802),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net802),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net802),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(rst_n),
    .X(net803));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(tmds_b));
 sg13g2_buf_1 output4 (.A(net4),
    .X(tmds_clk));
 sg13g2_buf_1 output5 (.A(net5),
    .X(tmds_g));
 sg13g2_buf_1 output6 (.A(net6),
    .X(tmds_r));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[7]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_bagel_21 (.L_LO(net21));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_3_0__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_3_4__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_1 clkload6 (.A(clknet_3_6__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\clockdiv.q2 ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0623_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold3 (.A(\serialize.n420[1] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold4 (.A(\serialize.n420[0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold5 (.A(\serialize.n420[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold6 (.A(\serialize.n420[3] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold7 (.A(\serialize.n420[4] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold8 (.A(\serialize.bit_cnt[0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold9 (.A(\serialize.n414[3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold10 (.A(\serialize.n420[6] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold11 (.A(\serialize.n431[6] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold12 (.A(\serialize.n414[1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold13 (.A(\serialize.n417[6] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold14 (.A(\serialize.n411[6] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold15 (.A(\serialize.n427[6] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold16 (.A(\serialize.n414[5] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold17 (.A(\serialize.n414[4] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold18 (.A(\serialize.n411[5] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold19 (.A(\serialize.n411[7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold20 (.A(\serialize.n414[0] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold21 (.A(\serialize.n417[1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold22 (.A(\serialize.n414[6] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold23 (.A(\serialize.n428[6] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold24 (.A(\serialize.bit_cnt[1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold25 (.A(\serialize.n410 ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold26 (.A(\serialize.n411[2] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold27 (.A(\serialize.n411[1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold28 (.A(\serialize.n417[0] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold29 (.A(\clockdiv.q0 ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold30 (.A(\serialize.n411[4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold31 (.A(\serialize.n417[3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold32 (.A(\serialize.n411[3] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold33 (.A(\serialize.n411[0] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold34 (.A(\serialize.n414[7] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold35 (.A(\serialize.n414[2] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold36 (.A(\serialize.n417[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold37 (.A(\serialize.n417[7] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold38 (.A(\serialize.n417[4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0004_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold40 (.A(\serialize.n417[5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0004_),
    .X(net446));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_44 ();
 sg13g2_fill_2 FILLER_0_53 ();
 sg13g2_fill_1 FILLER_0_55 ();
 sg13g2_decap_8 FILLER_0_60 ();
 sg13g2_decap_4 FILLER_0_67 ();
 sg13g2_fill_1 FILLER_0_71 ();
 sg13g2_fill_2 FILLER_0_77 ();
 sg13g2_fill_1 FILLER_0_79 ();
 sg13g2_decap_4 FILLER_0_85 ();
 sg13g2_fill_1 FILLER_0_89 ();
 sg13g2_decap_4 FILLER_0_95 ();
 sg13g2_fill_1 FILLER_0_99 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_fill_1 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_fill_1 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_156 ();
 sg13g2_decap_8 FILLER_0_163 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_fill_2 FILLER_0_198 ();
 sg13g2_fill_1 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_fill_1 FILLER_0_226 ();
 sg13g2_decap_4 FILLER_0_240 ();
 sg13g2_fill_1 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_4 FILLER_0_291 ();
 sg13g2_fill_2 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_343 ();
 sg13g2_fill_2 FILLER_0_372 ();
 sg13g2_fill_1 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_4 FILLER_0_386 ();
 sg13g2_fill_2 FILLER_0_390 ();
 sg13g2_fill_2 FILLER_0_396 ();
 sg13g2_fill_1 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_fill_2 FILLER_0_448 ();
 sg13g2_fill_1 FILLER_0_450 ();
 sg13g2_fill_1 FILLER_0_478 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_4 FILLER_0_525 ();
 sg13g2_fill_1 FILLER_0_529 ();
 sg13g2_decap_8 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_541 ();
 sg13g2_decap_8 FILLER_0_548 ();
 sg13g2_decap_8 FILLER_0_555 ();
 sg13g2_decap_8 FILLER_0_562 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_fill_2 FILLER_0_590 ();
 sg13g2_fill_1 FILLER_0_592 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_fill_2 FILLER_0_625 ();
 sg13g2_fill_1 FILLER_0_627 ();
 sg13g2_fill_2 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_8 FILLER_0_737 ();
 sg13g2_decap_8 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_751 ();
 sg13g2_decap_8 FILLER_0_758 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_8 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_779 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_884 ();
 sg13g2_decap_8 FILLER_0_891 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_905 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_8 FILLER_0_926 ();
 sg13g2_decap_8 FILLER_0_933 ();
 sg13g2_decap_8 FILLER_0_940 ();
 sg13g2_decap_8 FILLER_0_947 ();
 sg13g2_decap_8 FILLER_0_954 ();
 sg13g2_decap_8 FILLER_0_961 ();
 sg13g2_decap_8 FILLER_0_968 ();
 sg13g2_decap_8 FILLER_0_975 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_4 FILLER_0_1024 ();
 sg13g2_fill_1 FILLER_0_1028 ();
 sg13g2_decap_4 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_4 ();
 sg13g2_fill_1 FILLER_1_66 ();
 sg13g2_decap_4 FILLER_1_82 ();
 sg13g2_fill_2 FILLER_1_120 ();
 sg13g2_fill_1 FILLER_1_122 ();
 sg13g2_decap_4 FILLER_1_156 ();
 sg13g2_fill_2 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_169 ();
 sg13g2_fill_1 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_fill_2 FILLER_1_194 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_290 ();
 sg13g2_decap_4 FILLER_1_345 ();
 sg13g2_fill_1 FILLER_1_349 ();
 sg13g2_fill_2 FILLER_1_354 ();
 sg13g2_fill_1 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_446 ();
 sg13g2_fill_2 FILLER_1_453 ();
 sg13g2_fill_1 FILLER_1_455 ();
 sg13g2_decap_4 FILLER_1_460 ();
 sg13g2_fill_2 FILLER_1_495 ();
 sg13g2_fill_1 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_fill_1 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_662 ();
 sg13g2_decap_8 FILLER_1_669 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_4 FILLER_1_683 ();
 sg13g2_fill_2 FILLER_1_687 ();
 sg13g2_fill_1 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_8 FILLER_1_720 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_755 ();
 sg13g2_decap_8 FILLER_1_762 ();
 sg13g2_decap_8 FILLER_1_769 ();
 sg13g2_decap_8 FILLER_1_776 ();
 sg13g2_decap_8 FILLER_1_783 ();
 sg13g2_decap_8 FILLER_1_790 ();
 sg13g2_decap_8 FILLER_1_797 ();
 sg13g2_decap_8 FILLER_1_804 ();
 sg13g2_decap_8 FILLER_1_811 ();
 sg13g2_decap_8 FILLER_1_818 ();
 sg13g2_decap_8 FILLER_1_825 ();
 sg13g2_decap_8 FILLER_1_832 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_decap_8 FILLER_1_930 ();
 sg13g2_decap_8 FILLER_1_937 ();
 sg13g2_decap_8 FILLER_1_944 ();
 sg13g2_decap_8 FILLER_1_951 ();
 sg13g2_decap_8 FILLER_1_958 ();
 sg13g2_decap_8 FILLER_1_965 ();
 sg13g2_decap_8 FILLER_1_972 ();
 sg13g2_decap_8 FILLER_1_979 ();
 sg13g2_decap_8 FILLER_1_986 ();
 sg13g2_decap_8 FILLER_1_993 ();
 sg13g2_decap_8 FILLER_1_1000 ();
 sg13g2_decap_8 FILLER_1_1007 ();
 sg13g2_decap_8 FILLER_1_1014 ();
 sg13g2_decap_8 FILLER_1_1021 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_4 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_67 ();
 sg13g2_decap_4 FILLER_2_87 ();
 sg13g2_decap_4 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_103 ();
 sg13g2_decap_8 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_122 ();
 sg13g2_decap_8 FILLER_2_132 ();
 sg13g2_decap_8 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_146 ();
 sg13g2_decap_4 FILLER_2_153 ();
 sg13g2_decap_8 FILLER_2_185 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_fill_1 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_204 ();
 sg13g2_fill_1 FILLER_2_211 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_4 FILLER_2_279 ();
 sg13g2_fill_2 FILLER_2_283 ();
 sg13g2_decap_4 FILLER_2_289 ();
 sg13g2_fill_2 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_fill_1 FILLER_2_301 ();
 sg13g2_fill_2 FILLER_2_306 ();
 sg13g2_fill_1 FILLER_2_308 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_decap_4 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_4 FILLER_2_377 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_4 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_4 FILLER_2_414 ();
 sg13g2_fill_1 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_2_433 ();
 sg13g2_decap_4 FILLER_2_440 ();
 sg13g2_decap_8 FILLER_2_464 ();
 sg13g2_fill_2 FILLER_2_471 ();
 sg13g2_decap_8 FILLER_2_481 ();
 sg13g2_decap_8 FILLER_2_488 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_fill_2 FILLER_2_532 ();
 sg13g2_fill_1 FILLER_2_538 ();
 sg13g2_fill_2 FILLER_2_547 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_4 FILLER_2_564 ();
 sg13g2_fill_2 FILLER_2_568 ();
 sg13g2_decap_4 FILLER_2_578 ();
 sg13g2_fill_2 FILLER_2_582 ();
 sg13g2_decap_4 FILLER_2_610 ();
 sg13g2_fill_2 FILLER_2_622 ();
 sg13g2_fill_1 FILLER_2_624 ();
 sg13g2_fill_1 FILLER_2_641 ();
 sg13g2_fill_2 FILLER_2_650 ();
 sg13g2_fill_1 FILLER_2_652 ();
 sg13g2_decap_4 FILLER_2_681 ();
 sg13g2_fill_1 FILLER_2_702 ();
 sg13g2_decap_8 FILLER_2_716 ();
 sg13g2_decap_4 FILLER_2_723 ();
 sg13g2_fill_1 FILLER_2_727 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_8 FILLER_2_751 ();
 sg13g2_decap_8 FILLER_2_758 ();
 sg13g2_fill_2 FILLER_2_765 ();
 sg13g2_fill_2 FILLER_2_775 ();
 sg13g2_fill_1 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_787 ();
 sg13g2_decap_8 FILLER_2_794 ();
 sg13g2_decap_8 FILLER_2_801 ();
 sg13g2_fill_2 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_825 ();
 sg13g2_decap_8 FILLER_2_832 ();
 sg13g2_decap_8 FILLER_2_839 ();
 sg13g2_decap_8 FILLER_2_846 ();
 sg13g2_decap_8 FILLER_2_853 ();
 sg13g2_decap_8 FILLER_2_860 ();
 sg13g2_decap_8 FILLER_2_867 ();
 sg13g2_decap_8 FILLER_2_874 ();
 sg13g2_decap_8 FILLER_2_881 ();
 sg13g2_decap_8 FILLER_2_888 ();
 sg13g2_decap_8 FILLER_2_895 ();
 sg13g2_decap_8 FILLER_2_902 ();
 sg13g2_decap_8 FILLER_2_909 ();
 sg13g2_decap_8 FILLER_2_916 ();
 sg13g2_decap_8 FILLER_2_923 ();
 sg13g2_decap_8 FILLER_2_930 ();
 sg13g2_decap_8 FILLER_2_937 ();
 sg13g2_decap_8 FILLER_2_944 ();
 sg13g2_decap_8 FILLER_2_951 ();
 sg13g2_decap_8 FILLER_2_958 ();
 sg13g2_decap_8 FILLER_2_965 ();
 sg13g2_decap_8 FILLER_2_972 ();
 sg13g2_decap_8 FILLER_2_979 ();
 sg13g2_decap_8 FILLER_2_986 ();
 sg13g2_decap_8 FILLER_2_993 ();
 sg13g2_decap_8 FILLER_2_1000 ();
 sg13g2_decap_8 FILLER_2_1007 ();
 sg13g2_decap_8 FILLER_2_1014 ();
 sg13g2_decap_8 FILLER_2_1021 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_fill_1 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_20 ();
 sg13g2_decap_8 FILLER_3_27 ();
 sg13g2_fill_2 FILLER_3_34 ();
 sg13g2_fill_1 FILLER_3_36 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_56 ();
 sg13g2_fill_2 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_90 ();
 sg13g2_decap_8 FILLER_3_97 ();
 sg13g2_fill_1 FILLER_3_104 ();
 sg13g2_fill_2 FILLER_3_115 ();
 sg13g2_fill_1 FILLER_3_117 ();
 sg13g2_decap_4 FILLER_3_122 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_170 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_decap_4 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_222 ();
 sg13g2_fill_2 FILLER_3_238 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_279 ();
 sg13g2_decap_4 FILLER_3_307 ();
 sg13g2_fill_2 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_fill_2 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_fill_1 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_fill_1 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_446 ();
 sg13g2_decap_8 FILLER_3_453 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_4 FILLER_3_494 ();
 sg13g2_fill_1 FILLER_3_498 ();
 sg13g2_fill_1 FILLER_3_502 ();
 sg13g2_decap_8 FILLER_3_516 ();
 sg13g2_decap_8 FILLER_3_523 ();
 sg13g2_fill_2 FILLER_3_530 ();
 sg13g2_fill_1 FILLER_3_532 ();
 sg13g2_decap_4 FILLER_3_537 ();
 sg13g2_fill_1 FILLER_3_541 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_607 ();
 sg13g2_decap_8 FILLER_3_614 ();
 sg13g2_decap_8 FILLER_3_621 ();
 sg13g2_fill_2 FILLER_3_628 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_fill_1 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_656 ();
 sg13g2_decap_8 FILLER_3_663 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_decap_8 FILLER_3_677 ();
 sg13g2_decap_8 FILLER_3_684 ();
 sg13g2_fill_1 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_716 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_fill_2 FILLER_3_730 ();
 sg13g2_fill_1 FILLER_3_740 ();
 sg13g2_fill_1 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_decap_8 FILLER_3_841 ();
 sg13g2_decap_4 FILLER_3_848 ();
 sg13g2_fill_1 FILLER_3_852 ();
 sg13g2_decap_8 FILLER_3_862 ();
 sg13g2_decap_8 FILLER_3_869 ();
 sg13g2_decap_8 FILLER_3_876 ();
 sg13g2_decap_8 FILLER_3_883 ();
 sg13g2_decap_8 FILLER_3_890 ();
 sg13g2_decap_8 FILLER_3_897 ();
 sg13g2_decap_8 FILLER_3_904 ();
 sg13g2_decap_8 FILLER_3_911 ();
 sg13g2_decap_8 FILLER_3_918 ();
 sg13g2_decap_8 FILLER_3_925 ();
 sg13g2_decap_8 FILLER_3_932 ();
 sg13g2_decap_8 FILLER_3_939 ();
 sg13g2_decap_8 FILLER_3_946 ();
 sg13g2_decap_8 FILLER_3_953 ();
 sg13g2_decap_8 FILLER_3_960 ();
 sg13g2_decap_8 FILLER_3_967 ();
 sg13g2_decap_8 FILLER_3_974 ();
 sg13g2_decap_8 FILLER_3_981 ();
 sg13g2_decap_8 FILLER_3_988 ();
 sg13g2_decap_8 FILLER_3_995 ();
 sg13g2_decap_8 FILLER_3_1002 ();
 sg13g2_decap_8 FILLER_3_1009 ();
 sg13g2_decap_8 FILLER_3_1016 ();
 sg13g2_decap_4 FILLER_3_1023 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_decap_8 FILLER_4_31 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_decap_4 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_74 ();
 sg13g2_decap_4 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_160 ();
 sg13g2_decap_4 FILLER_4_172 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_181 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_decap_8 FILLER_4_195 ();
 sg13g2_decap_8 FILLER_4_202 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_decap_4 FILLER_4_228 ();
 sg13g2_fill_2 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_fill_1 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_4 FILLER_4_299 ();
 sg13g2_fill_2 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_311 ();
 sg13g2_decap_4 FILLER_4_333 ();
 sg13g2_fill_2 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_fill_1 FILLER_4_404 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_4 FILLER_4_423 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_decap_4 FILLER_4_470 ();
 sg13g2_fill_1 FILLER_4_474 ();
 sg13g2_decap_8 FILLER_4_506 ();
 sg13g2_fill_2 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_565 ();
 sg13g2_decap_8 FILLER_4_572 ();
 sg13g2_decap_4 FILLER_4_579 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_fill_2 FILLER_4_623 ();
 sg13g2_decap_4 FILLER_4_630 ();
 sg13g2_fill_2 FILLER_4_644 ();
 sg13g2_fill_1 FILLER_4_646 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_decap_4 FILLER_4_682 ();
 sg13g2_fill_1 FILLER_4_690 ();
 sg13g2_fill_2 FILLER_4_699 ();
 sg13g2_fill_1 FILLER_4_701 ();
 sg13g2_decap_8 FILLER_4_715 ();
 sg13g2_decap_8 FILLER_4_722 ();
 sg13g2_decap_8 FILLER_4_729 ();
 sg13g2_decap_4 FILLER_4_736 ();
 sg13g2_fill_2 FILLER_4_744 ();
 sg13g2_fill_2 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_793 ();
 sg13g2_fill_1 FILLER_4_800 ();
 sg13g2_decap_4 FILLER_4_825 ();
 sg13g2_decap_4 FILLER_4_850 ();
 sg13g2_decap_8 FILLER_4_880 ();
 sg13g2_decap_8 FILLER_4_887 ();
 sg13g2_decap_8 FILLER_4_894 ();
 sg13g2_decap_8 FILLER_4_901 ();
 sg13g2_decap_8 FILLER_4_908 ();
 sg13g2_decap_8 FILLER_4_915 ();
 sg13g2_decap_8 FILLER_4_922 ();
 sg13g2_decap_8 FILLER_4_929 ();
 sg13g2_decap_8 FILLER_4_936 ();
 sg13g2_decap_8 FILLER_4_943 ();
 sg13g2_decap_8 FILLER_4_950 ();
 sg13g2_decap_8 FILLER_4_957 ();
 sg13g2_decap_8 FILLER_4_964 ();
 sg13g2_decap_8 FILLER_4_971 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_8 FILLER_4_992 ();
 sg13g2_decap_8 FILLER_4_999 ();
 sg13g2_decap_8 FILLER_4_1006 ();
 sg13g2_decap_8 FILLER_4_1013 ();
 sg13g2_decap_8 FILLER_4_1020 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_fill_2 FILLER_5_8 ();
 sg13g2_fill_1 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_19 ();
 sg13g2_fill_2 FILLER_5_26 ();
 sg13g2_decap_8 FILLER_5_38 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_2 FILLER_5_79 ();
 sg13g2_fill_2 FILLER_5_85 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_decap_4 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_decap_8 FILLER_5_101 ();
 sg13g2_fill_2 FILLER_5_108 ();
 sg13g2_fill_1 FILLER_5_110 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_decap_4 FILLER_5_129 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_decap_4 FILLER_5_146 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_decap_4 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_fill_1 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_4 FILLER_5_366 ();
 sg13g2_fill_1 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_fill_1 FILLER_5_433 ();
 sg13g2_fill_2 FILLER_5_438 ();
 sg13g2_fill_1 FILLER_5_440 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_4 FILLER_5_466 ();
 sg13g2_fill_2 FILLER_5_470 ();
 sg13g2_fill_2 FILLER_5_482 ();
 sg13g2_decap_8 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_495 ();
 sg13g2_decap_8 FILLER_5_502 ();
 sg13g2_fill_2 FILLER_5_509 ();
 sg13g2_fill_1 FILLER_5_511 ();
 sg13g2_fill_2 FILLER_5_516 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_fill_2 FILLER_5_536 ();
 sg13g2_fill_2 FILLER_5_554 ();
 sg13g2_fill_1 FILLER_5_556 ();
 sg13g2_fill_2 FILLER_5_590 ();
 sg13g2_fill_1 FILLER_5_592 ();
 sg13g2_fill_1 FILLER_5_597 ();
 sg13g2_fill_1 FILLER_5_636 ();
 sg13g2_fill_2 FILLER_5_651 ();
 sg13g2_fill_1 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_679 ();
 sg13g2_fill_1 FILLER_5_685 ();
 sg13g2_fill_2 FILLER_5_699 ();
 sg13g2_decap_4 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_4 FILLER_5_756 ();
 sg13g2_fill_1 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_4 FILLER_5_777 ();
 sg13g2_fill_1 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_787 ();
 sg13g2_decap_8 FILLER_5_794 ();
 sg13g2_decap_4 FILLER_5_813 ();
 sg13g2_decap_4 FILLER_5_825 ();
 sg13g2_fill_1 FILLER_5_829 ();
 sg13g2_decap_8 FILLER_5_853 ();
 sg13g2_decap_8 FILLER_5_883 ();
 sg13g2_decap_8 FILLER_5_890 ();
 sg13g2_decap_8 FILLER_5_897 ();
 sg13g2_decap_8 FILLER_5_904 ();
 sg13g2_decap_8 FILLER_5_911 ();
 sg13g2_decap_8 FILLER_5_918 ();
 sg13g2_decap_8 FILLER_5_925 ();
 sg13g2_decap_8 FILLER_5_932 ();
 sg13g2_decap_8 FILLER_5_939 ();
 sg13g2_decap_8 FILLER_5_946 ();
 sg13g2_decap_8 FILLER_5_953 ();
 sg13g2_decap_8 FILLER_5_960 ();
 sg13g2_decap_8 FILLER_5_967 ();
 sg13g2_decap_8 FILLER_5_974 ();
 sg13g2_decap_8 FILLER_5_981 ();
 sg13g2_decap_8 FILLER_5_988 ();
 sg13g2_decap_8 FILLER_5_995 ();
 sg13g2_decap_8 FILLER_5_1002 ();
 sg13g2_decap_8 FILLER_5_1009 ();
 sg13g2_decap_8 FILLER_5_1016 ();
 sg13g2_decap_4 FILLER_5_1023 ();
 sg13g2_fill_2 FILLER_5_1027 ();
 sg13g2_decap_8 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_decap_4 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_43 ();
 sg13g2_fill_2 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_fill_2 FILLER_6_66 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_106 ();
 sg13g2_decap_4 FILLER_6_113 ();
 sg13g2_fill_2 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_174 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_decap_4 FILLER_6_187 ();
 sg13g2_decap_4 FILLER_6_195 ();
 sg13g2_decap_4 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_4 FILLER_6_262 ();
 sg13g2_fill_2 FILLER_6_293 ();
 sg13g2_fill_1 FILLER_6_295 ();
 sg13g2_decap_4 FILLER_6_313 ();
 sg13g2_decap_4 FILLER_6_330 ();
 sg13g2_fill_2 FILLER_6_334 ();
 sg13g2_decap_4 FILLER_6_373 ();
 sg13g2_fill_2 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_fill_1 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_fill_2 FILLER_6_416 ();
 sg13g2_decap_4 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_426 ();
 sg13g2_fill_2 FILLER_6_437 ();
 sg13g2_decap_4 FILLER_6_449 ();
 sg13g2_fill_1 FILLER_6_453 ();
 sg13g2_decap_8 FILLER_6_458 ();
 sg13g2_decap_8 FILLER_6_465 ();
 sg13g2_decap_4 FILLER_6_472 ();
 sg13g2_decap_8 FILLER_6_489 ();
 sg13g2_fill_2 FILLER_6_519 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_fill_1 FILLER_6_532 ();
 sg13g2_decap_4 FILLER_6_542 ();
 sg13g2_decap_4 FILLER_6_554 ();
 sg13g2_fill_1 FILLER_6_558 ();
 sg13g2_decap_4 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_572 ();
 sg13g2_decap_8 FILLER_6_579 ();
 sg13g2_decap_8 FILLER_6_586 ();
 sg13g2_fill_2 FILLER_6_593 ();
 sg13g2_decap_4 FILLER_6_604 ();
 sg13g2_decap_8 FILLER_6_612 ();
 sg13g2_decap_8 FILLER_6_619 ();
 sg13g2_decap_8 FILLER_6_626 ();
 sg13g2_fill_1 FILLER_6_633 ();
 sg13g2_fill_2 FILLER_6_647 ();
 sg13g2_fill_1 FILLER_6_676 ();
 sg13g2_fill_2 FILLER_6_687 ();
 sg13g2_fill_1 FILLER_6_689 ();
 sg13g2_fill_1 FILLER_6_695 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_fill_1 FILLER_6_728 ();
 sg13g2_fill_1 FILLER_6_756 ();
 sg13g2_decap_4 FILLER_6_795 ();
 sg13g2_fill_1 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_856 ();
 sg13g2_decap_4 FILLER_6_863 ();
 sg13g2_fill_2 FILLER_6_867 ();
 sg13g2_fill_1 FILLER_6_887 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_4 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1023 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_10 ();
 sg13g2_fill_1 FILLER_7_12 ();
 sg13g2_decap_4 FILLER_7_17 ();
 sg13g2_decap_8 FILLER_7_75 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_120 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_decap_8 FILLER_7_163 ();
 sg13g2_decap_4 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_178 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_decap_4 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_4 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_4 FILLER_7_372 ();
 sg13g2_fill_2 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_fill_2 FILLER_7_440 ();
 sg13g2_fill_1 FILLER_7_442 ();
 sg13g2_decap_4 FILLER_7_470 ();
 sg13g2_fill_2 FILLER_7_474 ();
 sg13g2_fill_2 FILLER_7_503 ();
 sg13g2_fill_1 FILLER_7_505 ();
 sg13g2_fill_2 FILLER_7_533 ();
 sg13g2_fill_1 FILLER_7_535 ();
 sg13g2_fill_2 FILLER_7_540 ();
 sg13g2_decap_8 FILLER_7_555 ();
 sg13g2_decap_8 FILLER_7_562 ();
 sg13g2_decap_8 FILLER_7_573 ();
 sg13g2_decap_8 FILLER_7_580 ();
 sg13g2_fill_2 FILLER_7_587 ();
 sg13g2_fill_1 FILLER_7_597 ();
 sg13g2_fill_2 FILLER_7_610 ();
 sg13g2_fill_1 FILLER_7_612 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_fill_2 FILLER_7_665 ();
 sg13g2_decap_4 FILLER_7_692 ();
 sg13g2_fill_2 FILLER_7_696 ();
 sg13g2_fill_2 FILLER_7_702 ();
 sg13g2_decap_8 FILLER_7_709 ();
 sg13g2_decap_8 FILLER_7_716 ();
 sg13g2_decap_4 FILLER_7_723 ();
 sg13g2_decap_8 FILLER_7_752 ();
 sg13g2_decap_4 FILLER_7_759 ();
 sg13g2_decap_8 FILLER_7_781 ();
 sg13g2_decap_8 FILLER_7_788 ();
 sg13g2_fill_2 FILLER_7_795 ();
 sg13g2_fill_1 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_4 FILLER_7_826 ();
 sg13g2_fill_1 FILLER_7_830 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_fill_2 FILLER_7_859 ();
 sg13g2_decap_4 FILLER_7_866 ();
 sg13g2_fill_2 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_decap_8 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_decap_8 FILLER_7_954 ();
 sg13g2_decap_8 FILLER_7_961 ();
 sg13g2_decap_8 FILLER_7_968 ();
 sg13g2_decap_8 FILLER_7_975 ();
 sg13g2_decap_8 FILLER_7_982 ();
 sg13g2_decap_8 FILLER_7_989 ();
 sg13g2_decap_8 FILLER_7_996 ();
 sg13g2_decap_8 FILLER_7_1003 ();
 sg13g2_decap_8 FILLER_7_1010 ();
 sg13g2_decap_8 FILLER_7_1017 ();
 sg13g2_decap_4 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_4 FILLER_8_11 ();
 sg13g2_fill_1 FILLER_8_15 ();
 sg13g2_decap_4 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_24 ();
 sg13g2_decap_4 FILLER_8_39 ();
 sg13g2_fill_1 FILLER_8_43 ();
 sg13g2_decap_8 FILLER_8_66 ();
 sg13g2_fill_2 FILLER_8_73 ();
 sg13g2_decap_4 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_83 ();
 sg13g2_fill_1 FILLER_8_89 ();
 sg13g2_decap_4 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_138 ();
 sg13g2_decap_8 FILLER_8_145 ();
 sg13g2_decap_4 FILLER_8_152 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_decap_4 FILLER_8_205 ();
 sg13g2_fill_2 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_decap_4 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_4 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_2 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_fill_2 FILLER_8_429 ();
 sg13g2_fill_1 FILLER_8_431 ();
 sg13g2_fill_2 FILLER_8_436 ();
 sg13g2_fill_1 FILLER_8_438 ();
 sg13g2_decap_4 FILLER_8_443 ();
 sg13g2_fill_1 FILLER_8_447 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_4 FILLER_8_459 ();
 sg13g2_fill_1 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_478 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_489 ();
 sg13g2_decap_8 FILLER_8_496 ();
 sg13g2_decap_4 FILLER_8_503 ();
 sg13g2_fill_2 FILLER_8_515 ();
 sg13g2_fill_1 FILLER_8_517 ();
 sg13g2_fill_1 FILLER_8_531 ();
 sg13g2_decap_4 FILLER_8_560 ();
 sg13g2_fill_1 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_604 ();
 sg13g2_fill_2 FILLER_8_627 ();
 sg13g2_fill_1 FILLER_8_629 ();
 sg13g2_fill_2 FILLER_8_637 ();
 sg13g2_fill_1 FILLER_8_639 ();
 sg13g2_decap_8 FILLER_8_650 ();
 sg13g2_decap_8 FILLER_8_657 ();
 sg13g2_decap_8 FILLER_8_664 ();
 sg13g2_fill_2 FILLER_8_671 ();
 sg13g2_decap_8 FILLER_8_684 ();
 sg13g2_decap_8 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_715 ();
 sg13g2_fill_2 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_751 ();
 sg13g2_decap_4 FILLER_8_758 ();
 sg13g2_fill_2 FILLER_8_762 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_4 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_820 ();
 sg13g2_decap_4 FILLER_8_827 ();
 sg13g2_fill_1 FILLER_8_831 ();
 sg13g2_decap_4 FILLER_8_848 ();
 sg13g2_fill_2 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_870 ();
 sg13g2_decap_8 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_891 ();
 sg13g2_decap_8 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_905 ();
 sg13g2_decap_8 FILLER_8_912 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_decap_8 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_933 ();
 sg13g2_decap_8 FILLER_8_940 ();
 sg13g2_decap_8 FILLER_8_947 ();
 sg13g2_decap_8 FILLER_8_954 ();
 sg13g2_decap_8 FILLER_8_961 ();
 sg13g2_decap_8 FILLER_8_968 ();
 sg13g2_decap_8 FILLER_8_975 ();
 sg13g2_decap_8 FILLER_8_982 ();
 sg13g2_decap_8 FILLER_8_989 ();
 sg13g2_decap_8 FILLER_8_996 ();
 sg13g2_decap_8 FILLER_8_1003 ();
 sg13g2_decap_8 FILLER_8_1010 ();
 sg13g2_decap_8 FILLER_8_1017 ();
 sg13g2_decap_4 FILLER_8_1024 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_43 ();
 sg13g2_decap_8 FILLER_9_50 ();
 sg13g2_decap_8 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_64 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_2 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_93 ();
 sg13g2_decap_8 FILLER_9_121 ();
 sg13g2_decap_4 FILLER_9_128 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_4 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_187 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_201 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_4 FILLER_9_249 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_2 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_4 FILLER_9_301 ();
 sg13g2_fill_2 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_342 ();
 sg13g2_decap_4 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_fill_2 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_fill_2 FILLER_9_434 ();
 sg13g2_fill_1 FILLER_9_436 ();
 sg13g2_decap_4 FILLER_9_452 ();
 sg13g2_fill_1 FILLER_9_456 ();
 sg13g2_fill_2 FILLER_9_492 ();
 sg13g2_decap_8 FILLER_9_498 ();
 sg13g2_decap_8 FILLER_9_505 ();
 sg13g2_decap_8 FILLER_9_512 ();
 sg13g2_decap_8 FILLER_9_519 ();
 sg13g2_fill_2 FILLER_9_526 ();
 sg13g2_fill_2 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_fill_2 FILLER_9_567 ();
 sg13g2_fill_1 FILLER_9_569 ();
 sg13g2_decap_4 FILLER_9_574 ();
 sg13g2_fill_1 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_fill_2 FILLER_9_631 ();
 sg13g2_fill_1 FILLER_9_633 ();
 sg13g2_fill_2 FILLER_9_667 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_fill_1 FILLER_9_740 ();
 sg13g2_decap_8 FILLER_9_748 ();
 sg13g2_fill_2 FILLER_9_755 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_4 FILLER_9_795 ();
 sg13g2_fill_1 FILLER_9_799 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_4 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_848 ();
 sg13g2_decap_4 FILLER_9_855 ();
 sg13g2_fill_2 FILLER_9_859 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_fill_2 FILLER_9_889 ();
 sg13g2_fill_1 FILLER_9_891 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_10_16 ();
 sg13g2_decap_8 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_30 ();
 sg13g2_decap_8 FILLER_10_51 ();
 sg13g2_decap_4 FILLER_10_58 ();
 sg13g2_decap_4 FILLER_10_94 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_4 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_decap_4 FILLER_10_230 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_281 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_1 FILLER_10_372 ();
 sg13g2_fill_2 FILLER_10_377 ();
 sg13g2_decap_4 FILLER_10_389 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_decap_4 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_426 ();
 sg13g2_decap_4 FILLER_10_454 ();
 sg13g2_fill_1 FILLER_10_458 ();
 sg13g2_decap_8 FILLER_10_463 ();
 sg13g2_fill_1 FILLER_10_470 ();
 sg13g2_fill_1 FILLER_10_476 ();
 sg13g2_fill_2 FILLER_10_487 ();
 sg13g2_decap_4 FILLER_10_521 ();
 sg13g2_fill_2 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_559 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_decap_4 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_fill_1 FILLER_10_631 ();
 sg13g2_decap_8 FILLER_10_646 ();
 sg13g2_decap_8 FILLER_10_653 ();
 sg13g2_decap_4 FILLER_10_660 ();
 sg13g2_decap_4 FILLER_10_682 ();
 sg13g2_fill_2 FILLER_10_686 ();
 sg13g2_decap_4 FILLER_10_701 ();
 sg13g2_decap_4 FILLER_10_713 ();
 sg13g2_decap_8 FILLER_10_726 ();
 sg13g2_fill_1 FILLER_10_733 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_4 FILLER_10_756 ();
 sg13g2_fill_1 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_fill_2 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_4 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_fill_2 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_856 ();
 sg13g2_fill_2 FILLER_10_879 ();
 sg13g2_fill_1 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_905 ();
 sg13g2_decap_8 FILLER_10_912 ();
 sg13g2_decap_8 FILLER_10_919 ();
 sg13g2_decap_8 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_933 ();
 sg13g2_decap_8 FILLER_10_940 ();
 sg13g2_decap_8 FILLER_10_947 ();
 sg13g2_decap_8 FILLER_10_954 ();
 sg13g2_decap_8 FILLER_10_961 ();
 sg13g2_decap_8 FILLER_10_968 ();
 sg13g2_decap_8 FILLER_10_975 ();
 sg13g2_decap_8 FILLER_10_982 ();
 sg13g2_decap_8 FILLER_10_989 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_8 FILLER_10_1003 ();
 sg13g2_decap_8 FILLER_10_1010 ();
 sg13g2_decap_8 FILLER_10_1017 ();
 sg13g2_decap_4 FILLER_10_1024 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_fill_2 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_4 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_127 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_decap_4 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_decap_4 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_4 FILLER_11_310 ();
 sg13g2_fill_2 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_4 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_4 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_386 ();
 sg13g2_decap_4 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_11_415 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_4 FILLER_11_452 ();
 sg13g2_decap_4 FILLER_11_493 ();
 sg13g2_fill_2 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_503 ();
 sg13g2_decap_8 FILLER_11_510 ();
 sg13g2_decap_8 FILLER_11_517 ();
 sg13g2_decap_8 FILLER_11_524 ();
 sg13g2_fill_1 FILLER_11_531 ();
 sg13g2_fill_1 FILLER_11_540 ();
 sg13g2_decap_8 FILLER_11_551 ();
 sg13g2_decap_4 FILLER_11_558 ();
 sg13g2_decap_4 FILLER_11_603 ();
 sg13g2_fill_2 FILLER_11_623 ();
 sg13g2_fill_1 FILLER_11_625 ();
 sg13g2_decap_4 FILLER_11_631 ();
 sg13g2_fill_1 FILLER_11_635 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_4 FILLER_11_654 ();
 sg13g2_decap_4 FILLER_11_662 ();
 sg13g2_fill_1 FILLER_11_666 ();
 sg13g2_fill_2 FILLER_11_679 ();
 sg13g2_fill_1 FILLER_11_681 ();
 sg13g2_fill_2 FILLER_11_692 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_decap_4 FILLER_11_709 ();
 sg13g2_decap_4 FILLER_11_716 ();
 sg13g2_fill_2 FILLER_11_720 ();
 sg13g2_fill_2 FILLER_11_728 ();
 sg13g2_fill_1 FILLER_11_730 ();
 sg13g2_fill_1 FILLER_11_744 ();
 sg13g2_decap_8 FILLER_11_751 ();
 sg13g2_decap_4 FILLER_11_758 ();
 sg13g2_fill_2 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_778 ();
 sg13g2_decap_8 FILLER_11_785 ();
 sg13g2_decap_8 FILLER_11_792 ();
 sg13g2_decap_4 FILLER_11_799 ();
 sg13g2_fill_2 FILLER_11_819 ();
 sg13g2_fill_1 FILLER_11_821 ();
 sg13g2_decap_4 FILLER_11_847 ();
 sg13g2_fill_2 FILLER_11_851 ();
 sg13g2_decap_4 FILLER_11_881 ();
 sg13g2_fill_2 FILLER_11_885 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_9 ();
 sg13g2_decap_8 FILLER_12_16 ();
 sg13g2_decap_8 FILLER_12_23 ();
 sg13g2_decap_8 FILLER_12_30 ();
 sg13g2_decap_4 FILLER_12_37 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_57 ();
 sg13g2_fill_2 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_66 ();
 sg13g2_decap_4 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_decap_4 FILLER_12_90 ();
 sg13g2_decap_4 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_decap_8 FILLER_12_114 ();
 sg13g2_decap_8 FILLER_12_121 ();
 sg13g2_decap_4 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_decap_4 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_4 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_fill_2 FILLER_12_306 ();
 sg13g2_decap_4 FILLER_12_333 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_2 FILLER_12_392 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_4 FILLER_12_414 ();
 sg13g2_fill_1 FILLER_12_418 ();
 sg13g2_fill_2 FILLER_12_425 ();
 sg13g2_decap_8 FILLER_12_432 ();
 sg13g2_fill_2 FILLER_12_439 ();
 sg13g2_fill_1 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_fill_2 FILLER_12_459 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_decap_4 FILLER_12_466 ();
 sg13g2_fill_1 FILLER_12_470 ();
 sg13g2_fill_2 FILLER_12_475 ();
 sg13g2_fill_1 FILLER_12_477 ();
 sg13g2_decap_8 FILLER_12_482 ();
 sg13g2_decap_4 FILLER_12_489 ();
 sg13g2_fill_1 FILLER_12_493 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_4 FILLER_12_529 ();
 sg13g2_fill_1 FILLER_12_538 ();
 sg13g2_decap_8 FILLER_12_570 ();
 sg13g2_decap_8 FILLER_12_577 ();
 sg13g2_decap_8 FILLER_12_594 ();
 sg13g2_decap_8 FILLER_12_601 ();
 sg13g2_decap_4 FILLER_12_608 ();
 sg13g2_decap_8 FILLER_12_624 ();
 sg13g2_decap_8 FILLER_12_631 ();
 sg13g2_fill_1 FILLER_12_638 ();
 sg13g2_decap_8 FILLER_12_681 ();
 sg13g2_decap_4 FILLER_12_688 ();
 sg13g2_decap_4 FILLER_12_696 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_decap_4 FILLER_12_719 ();
 sg13g2_fill_1 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_786 ();
 sg13g2_decap_8 FILLER_12_793 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_fill_2 FILLER_12_828 ();
 sg13g2_fill_1 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_fill_2 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_873 ();
 sg13g2_decap_8 FILLER_12_880 ();
 sg13g2_decap_8 FILLER_12_911 ();
 sg13g2_decap_8 FILLER_12_918 ();
 sg13g2_decap_8 FILLER_12_925 ();
 sg13g2_decap_8 FILLER_12_932 ();
 sg13g2_decap_8 FILLER_12_939 ();
 sg13g2_decap_8 FILLER_12_946 ();
 sg13g2_decap_8 FILLER_12_953 ();
 sg13g2_decap_8 FILLER_12_960 ();
 sg13g2_decap_8 FILLER_12_967 ();
 sg13g2_decap_8 FILLER_12_974 ();
 sg13g2_decap_8 FILLER_12_981 ();
 sg13g2_decap_8 FILLER_12_988 ();
 sg13g2_decap_8 FILLER_12_995 ();
 sg13g2_decap_8 FILLER_12_1002 ();
 sg13g2_decap_8 FILLER_12_1009 ();
 sg13g2_decap_8 FILLER_12_1016 ();
 sg13g2_decap_4 FILLER_12_1023 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_decap_4 FILLER_13_8 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_fill_2 FILLER_13_136 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_decap_4 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_decap_4 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_fill_1 FILLER_13_420 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_443 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_fill_2 FILLER_13_483 ();
 sg13g2_fill_2 FILLER_13_489 ();
 sg13g2_fill_1 FILLER_13_496 ();
 sg13g2_decap_8 FILLER_13_505 ();
 sg13g2_fill_2 FILLER_13_512 ();
 sg13g2_decap_4 FILLER_13_520 ();
 sg13g2_decap_8 FILLER_13_557 ();
 sg13g2_decap_8 FILLER_13_564 ();
 sg13g2_fill_2 FILLER_13_571 ();
 sg13g2_fill_1 FILLER_13_573 ();
 sg13g2_fill_2 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_619 ();
 sg13g2_fill_2 FILLER_13_626 ();
 sg13g2_fill_1 FILLER_13_628 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_fill_2 FILLER_13_656 ();
 sg13g2_fill_1 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_666 ();
 sg13g2_decap_8 FILLER_13_673 ();
 sg13g2_decap_4 FILLER_13_680 ();
 sg13g2_fill_2 FILLER_13_701 ();
 sg13g2_decap_8 FILLER_13_713 ();
 sg13g2_decap_8 FILLER_13_720 ();
 sg13g2_decap_4 FILLER_13_727 ();
 sg13g2_decap_8 FILLER_13_748 ();
 sg13g2_decap_8 FILLER_13_755 ();
 sg13g2_decap_8 FILLER_13_762 ();
 sg13g2_fill_2 FILLER_13_769 ();
 sg13g2_fill_1 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_4 FILLER_13_795 ();
 sg13g2_decap_4 FILLER_13_819 ();
 sg13g2_fill_1 FILLER_13_823 ();
 sg13g2_decap_4 FILLER_13_847 ();
 sg13g2_fill_1 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_877 ();
 sg13g2_decap_4 FILLER_13_884 ();
 sg13g2_fill_1 FILLER_13_888 ();
 sg13g2_decap_8 FILLER_13_916 ();
 sg13g2_decap_8 FILLER_13_923 ();
 sg13g2_decap_8 FILLER_13_930 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_8 FILLER_13_951 ();
 sg13g2_decap_8 FILLER_13_958 ();
 sg13g2_decap_8 FILLER_13_965 ();
 sg13g2_decap_8 FILLER_13_972 ();
 sg13g2_decap_8 FILLER_13_979 ();
 sg13g2_decap_8 FILLER_13_986 ();
 sg13g2_decap_8 FILLER_13_993 ();
 sg13g2_decap_8 FILLER_13_1000 ();
 sg13g2_decap_8 FILLER_13_1007 ();
 sg13g2_decap_8 FILLER_13_1014 ();
 sg13g2_decap_8 FILLER_13_1021 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_decap_8 FILLER_14_59 ();
 sg13g2_decap_8 FILLER_14_66 ();
 sg13g2_fill_1 FILLER_14_73 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_99 ();
 sg13g2_decap_4 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_fill_1 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_decap_4 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_4 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_4 FILLER_14_324 ();
 sg13g2_decap_4 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_342 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_4 FILLER_14_439 ();
 sg13g2_decap_8 FILLER_14_460 ();
 sg13g2_decap_8 FILLER_14_467 ();
 sg13g2_decap_4 FILLER_14_474 ();
 sg13g2_fill_1 FILLER_14_478 ();
 sg13g2_fill_2 FILLER_14_500 ();
 sg13g2_fill_2 FILLER_14_516 ();
 sg13g2_fill_1 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_fill_2 FILLER_14_532 ();
 sg13g2_fill_1 FILLER_14_534 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_fill_1 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_564 ();
 sg13g2_decap_8 FILLER_14_571 ();
 sg13g2_fill_1 FILLER_14_578 ();
 sg13g2_decap_4 FILLER_14_583 ();
 sg13g2_fill_2 FILLER_14_587 ();
 sg13g2_decap_8 FILLER_14_593 ();
 sg13g2_fill_1 FILLER_14_600 ();
 sg13g2_decap_4 FILLER_14_618 ();
 sg13g2_fill_2 FILLER_14_622 ();
 sg13g2_fill_2 FILLER_14_684 ();
 sg13g2_fill_1 FILLER_14_686 ();
 sg13g2_fill_1 FILLER_14_699 ();
 sg13g2_decap_4 FILLER_14_721 ();
 sg13g2_fill_2 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_750 ();
 sg13g2_decap_8 FILLER_14_757 ();
 sg13g2_fill_1 FILLER_14_764 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_800 ();
 sg13g2_fill_1 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_fill_2 FILLER_14_826 ();
 sg13g2_fill_1 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_4 FILLER_14_849 ();
 sg13g2_fill_1 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_fill_2 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_915 ();
 sg13g2_decap_8 FILLER_14_922 ();
 sg13g2_decap_8 FILLER_14_929 ();
 sg13g2_decap_8 FILLER_14_936 ();
 sg13g2_decap_8 FILLER_14_943 ();
 sg13g2_decap_8 FILLER_14_950 ();
 sg13g2_decap_8 FILLER_14_957 ();
 sg13g2_decap_8 FILLER_14_964 ();
 sg13g2_decap_8 FILLER_14_971 ();
 sg13g2_decap_8 FILLER_14_978 ();
 sg13g2_decap_8 FILLER_14_985 ();
 sg13g2_decap_8 FILLER_14_992 ();
 sg13g2_decap_8 FILLER_14_999 ();
 sg13g2_decap_8 FILLER_14_1006 ();
 sg13g2_decap_8 FILLER_14_1013 ();
 sg13g2_decap_8 FILLER_14_1020 ();
 sg13g2_fill_2 FILLER_14_1027 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_13 ();
 sg13g2_fill_2 FILLER_15_19 ();
 sg13g2_fill_1 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_decap_8 FILLER_15_31 ();
 sg13g2_decap_4 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_decap_4 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_decap_4 FILLER_15_160 ();
 sg13g2_decap_4 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_4 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_4 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_4 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_fill_2 FILLER_15_404 ();
 sg13g2_fill_2 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_15_435 ();
 sg13g2_decap_8 FILLER_15_442 ();
 sg13g2_decap_8 FILLER_15_449 ();
 sg13g2_fill_2 FILLER_15_456 ();
 sg13g2_fill_1 FILLER_15_458 ();
 sg13g2_fill_2 FILLER_15_487 ();
 sg13g2_fill_1 FILLER_15_489 ();
 sg13g2_fill_1 FILLER_15_518 ();
 sg13g2_fill_2 FILLER_15_546 ();
 sg13g2_fill_1 FILLER_15_548 ();
 sg13g2_fill_2 FILLER_15_553 ();
 sg13g2_fill_1 FILLER_15_555 ();
 sg13g2_decap_4 FILLER_15_562 ();
 sg13g2_fill_2 FILLER_15_566 ();
 sg13g2_decap_8 FILLER_15_580 ();
 sg13g2_decap_4 FILLER_15_587 ();
 sg13g2_fill_2 FILLER_15_591 ();
 sg13g2_fill_2 FILLER_15_597 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_fill_1 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_670 ();
 sg13g2_decap_8 FILLER_15_677 ();
 sg13g2_decap_4 FILLER_15_684 ();
 sg13g2_decap_8 FILLER_15_708 ();
 sg13g2_decap_4 FILLER_15_715 ();
 sg13g2_fill_1 FILLER_15_719 ();
 sg13g2_decap_4 FILLER_15_753 ();
 sg13g2_fill_2 FILLER_15_796 ();
 sg13g2_fill_1 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_4 FILLER_15_819 ();
 sg13g2_fill_1 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_fill_1 FILLER_15_856 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_938 ();
 sg13g2_decap_8 FILLER_15_945 ();
 sg13g2_decap_8 FILLER_15_952 ();
 sg13g2_decap_8 FILLER_15_959 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_decap_8 FILLER_15_973 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_8 FILLER_15_1001 ();
 sg13g2_decap_8 FILLER_15_1008 ();
 sg13g2_decap_8 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1022 ();
 sg13g2_decap_4 FILLER_16_27 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_39 ();
 sg13g2_decap_4 FILLER_16_51 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_148 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_4 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_decap_4 FILLER_16_314 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_430 ();
 sg13g2_fill_1 FILLER_16_432 ();
 sg13g2_fill_1 FILLER_16_443 ();
 sg13g2_fill_2 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_454 ();
 sg13g2_fill_1 FILLER_16_456 ();
 sg13g2_fill_1 FILLER_16_470 ();
 sg13g2_fill_2 FILLER_16_484 ();
 sg13g2_fill_1 FILLER_16_494 ();
 sg13g2_decap_4 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_503 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_fill_2 FILLER_16_536 ();
 sg13g2_fill_1 FILLER_16_538 ();
 sg13g2_fill_2 FILLER_16_627 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_decap_8 FILLER_16_666 ();
 sg13g2_decap_8 FILLER_16_673 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_fill_1 FILLER_16_738 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_4 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_789 ();
 sg13g2_decap_4 FILLER_16_796 ();
 sg13g2_fill_2 FILLER_16_800 ();
 sg13g2_fill_1 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_fill_1 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_fill_1 FILLER_16_850 ();
 sg13g2_decap_8 FILLER_16_874 ();
 sg13g2_decap_8 FILLER_16_881 ();
 sg13g2_fill_2 FILLER_16_888 ();
 sg13g2_fill_1 FILLER_16_890 ();
 sg13g2_decap_8 FILLER_16_922 ();
 sg13g2_decap_8 FILLER_16_929 ();
 sg13g2_decap_8 FILLER_16_936 ();
 sg13g2_decap_8 FILLER_16_943 ();
 sg13g2_decap_8 FILLER_16_950 ();
 sg13g2_decap_8 FILLER_16_957 ();
 sg13g2_decap_8 FILLER_16_964 ();
 sg13g2_decap_8 FILLER_16_971 ();
 sg13g2_decap_8 FILLER_16_978 ();
 sg13g2_decap_8 FILLER_16_985 ();
 sg13g2_decap_8 FILLER_16_992 ();
 sg13g2_decap_8 FILLER_16_999 ();
 sg13g2_decap_8 FILLER_16_1006 ();
 sg13g2_decap_8 FILLER_16_1013 ();
 sg13g2_decap_8 FILLER_16_1020 ();
 sg13g2_fill_2 FILLER_16_1027 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_9 ();
 sg13g2_decap_8 FILLER_17_16 ();
 sg13g2_fill_2 FILLER_17_23 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_17_66 ();
 sg13g2_decap_8 FILLER_17_71 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_4 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_433 ();
 sg13g2_fill_2 FILLER_17_437 ();
 sg13g2_decap_8 FILLER_17_470 ();
 sg13g2_decap_8 FILLER_17_477 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_fill_2 FILLER_17_535 ();
 sg13g2_fill_1 FILLER_17_537 ();
 sg13g2_decap_8 FILLER_17_551 ();
 sg13g2_decap_8 FILLER_17_558 ();
 sg13g2_decap_8 FILLER_17_565 ();
 sg13g2_decap_8 FILLER_17_590 ();
 sg13g2_decap_4 FILLER_17_597 ();
 sg13g2_fill_2 FILLER_17_607 ();
 sg13g2_decap_8 FILLER_17_622 ();
 sg13g2_fill_2 FILLER_17_629 ();
 sg13g2_fill_2 FILLER_17_644 ();
 sg13g2_fill_1 FILLER_17_646 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_fill_1 FILLER_17_689 ();
 sg13g2_fill_1 FILLER_17_695 ();
 sg13g2_fill_2 FILLER_17_701 ();
 sg13g2_fill_1 FILLER_17_703 ();
 sg13g2_decap_8 FILLER_17_709 ();
 sg13g2_decap_8 FILLER_17_716 ();
 sg13g2_decap_8 FILLER_17_723 ();
 sg13g2_fill_2 FILLER_17_751 ();
 sg13g2_fill_2 FILLER_17_767 ();
 sg13g2_fill_1 FILLER_17_769 ();
 sg13g2_decap_8 FILLER_17_789 ();
 sg13g2_fill_2 FILLER_17_796 ();
 sg13g2_fill_2 FILLER_17_820 ();
 sg13g2_fill_1 FILLER_17_822 ();
 sg13g2_fill_2 FILLER_17_841 ();
 sg13g2_fill_1 FILLER_17_860 ();
 sg13g2_decap_8 FILLER_17_883 ();
 sg13g2_decap_4 FILLER_17_890 ();
 sg13g2_fill_2 FILLER_17_894 ();
 sg13g2_decap_8 FILLER_17_921 ();
 sg13g2_decap_8 FILLER_17_928 ();
 sg13g2_decap_8 FILLER_17_935 ();
 sg13g2_decap_8 FILLER_17_942 ();
 sg13g2_decap_8 FILLER_17_949 ();
 sg13g2_decap_8 FILLER_17_956 ();
 sg13g2_decap_8 FILLER_17_963 ();
 sg13g2_decap_8 FILLER_17_970 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_984 ();
 sg13g2_decap_8 FILLER_17_991 ();
 sg13g2_decap_8 FILLER_17_998 ();
 sg13g2_decap_8 FILLER_17_1005 ();
 sg13g2_decap_8 FILLER_17_1012 ();
 sg13g2_decap_8 FILLER_17_1019 ();
 sg13g2_fill_2 FILLER_17_1026 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_decap_8 FILLER_18_8 ();
 sg13g2_decap_8 FILLER_18_15 ();
 sg13g2_fill_2 FILLER_18_22 ();
 sg13g2_fill_1 FILLER_18_24 ();
 sg13g2_decap_8 FILLER_18_45 ();
 sg13g2_decap_8 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_132 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_4 FILLER_18_258 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_4 FILLER_18_301 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_decap_4 FILLER_18_384 ();
 sg13g2_fill_2 FILLER_18_388 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_decap_4 FILLER_18_418 ();
 sg13g2_fill_2 FILLER_18_422 ();
 sg13g2_decap_8 FILLER_18_439 ();
 sg13g2_fill_2 FILLER_18_446 ();
 sg13g2_fill_1 FILLER_18_448 ();
 sg13g2_decap_4 FILLER_18_476 ();
 sg13g2_fill_2 FILLER_18_480 ();
 sg13g2_decap_4 FILLER_18_495 ();
 sg13g2_fill_2 FILLER_18_503 ();
 sg13g2_fill_1 FILLER_18_505 ();
 sg13g2_fill_2 FILLER_18_511 ();
 sg13g2_fill_1 FILLER_18_513 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_decap_8 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_4 FILLER_18_630 ();
 sg13g2_fill_1 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_640 ();
 sg13g2_fill_1 FILLER_18_642 ();
 sg13g2_fill_1 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_656 ();
 sg13g2_decap_8 FILLER_18_663 ();
 sg13g2_fill_2 FILLER_18_670 ();
 sg13g2_fill_2 FILLER_18_685 ();
 sg13g2_fill_1 FILLER_18_687 ();
 sg13g2_fill_1 FILLER_18_696 ();
 sg13g2_decap_4 FILLER_18_722 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_4 FILLER_18_766 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_fill_1 FILLER_18_795 ();
 sg13g2_fill_2 FILLER_18_809 ();
 sg13g2_decap_4 FILLER_18_823 ();
 sg13g2_fill_1 FILLER_18_827 ();
 sg13g2_decap_8 FILLER_18_832 ();
 sg13g2_decap_8 FILLER_18_839 ();
 sg13g2_decap_4 FILLER_18_846 ();
 sg13g2_decap_8 FILLER_18_876 ();
 sg13g2_decap_8 FILLER_18_883 ();
 sg13g2_decap_4 FILLER_18_890 ();
 sg13g2_decap_8 FILLER_18_917 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_decap_8 FILLER_18_938 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_decap_8 FILLER_18_952 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_10 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_19 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_4 FILLER_19_253 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_19_415 ();
 sg13g2_fill_2 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_439 ();
 sg13g2_fill_1 FILLER_19_443 ();
 sg13g2_fill_2 FILLER_19_471 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_fill_2 FILLER_19_533 ();
 sg13g2_fill_1 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_544 ();
 sg13g2_decap_8 FILLER_19_551 ();
 sg13g2_fill_1 FILLER_19_558 ();
 sg13g2_decap_4 FILLER_19_572 ();
 sg13g2_fill_1 FILLER_19_576 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_4 FILLER_19_595 ();
 sg13g2_fill_1 FILLER_19_615 ();
 sg13g2_fill_1 FILLER_19_631 ();
 sg13g2_decap_8 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_decap_4 FILLER_19_650 ();
 sg13g2_fill_1 FILLER_19_654 ();
 sg13g2_decap_8 FILLER_19_668 ();
 sg13g2_decap_8 FILLER_19_675 ();
 sg13g2_fill_1 FILLER_19_682 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_4 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_4 FILLER_19_763 ();
 sg13g2_fill_1 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_fill_2 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_815 ();
 sg13g2_fill_2 FILLER_19_822 ();
 sg13g2_fill_1 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_872 ();
 sg13g2_decap_8 FILLER_19_879 ();
 sg13g2_decap_4 FILLER_19_886 ();
 sg13g2_decap_8 FILLER_19_921 ();
 sg13g2_decap_8 FILLER_19_928 ();
 sg13g2_decap_8 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_942 ();
 sg13g2_decap_8 FILLER_19_949 ();
 sg13g2_decap_8 FILLER_19_956 ();
 sg13g2_decap_8 FILLER_19_963 ();
 sg13g2_decap_8 FILLER_19_970 ();
 sg13g2_decap_8 FILLER_19_977 ();
 sg13g2_decap_8 FILLER_19_984 ();
 sg13g2_decap_8 FILLER_19_991 ();
 sg13g2_decap_8 FILLER_19_998 ();
 sg13g2_decap_8 FILLER_19_1005 ();
 sg13g2_decap_8 FILLER_19_1012 ();
 sg13g2_decap_4 FILLER_19_1019 ();
 sg13g2_fill_2 FILLER_19_1023 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_38 ();
 sg13g2_fill_1 FILLER_20_43 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_decap_8 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_decap_4 FILLER_20_68 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_decap_8 FILLER_20_90 ();
 sg13g2_decap_8 FILLER_20_97 ();
 sg13g2_decap_4 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_decap_8 FILLER_20_122 ();
 sg13g2_decap_8 FILLER_20_129 ();
 sg13g2_decap_4 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_4 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_448 ();
 sg13g2_fill_2 FILLER_20_453 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_fill_2 FILLER_20_466 ();
 sg13g2_fill_1 FILLER_20_468 ();
 sg13g2_decap_8 FILLER_20_474 ();
 sg13g2_fill_2 FILLER_20_481 ();
 sg13g2_fill_1 FILLER_20_483 ();
 sg13g2_decap_4 FILLER_20_497 ();
 sg13g2_fill_1 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_507 ();
 sg13g2_decap_8 FILLER_20_514 ();
 sg13g2_decap_8 FILLER_20_521 ();
 sg13g2_decap_4 FILLER_20_528 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_decap_8 FILLER_20_573 ();
 sg13g2_decap_8 FILLER_20_580 ();
 sg13g2_decap_4 FILLER_20_587 ();
 sg13g2_decap_4 FILLER_20_608 ();
 sg13g2_fill_2 FILLER_20_612 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_4 FILLER_20_762 ();
 sg13g2_fill_1 FILLER_20_793 ();
 sg13g2_fill_1 FILLER_20_816 ();
 sg13g2_fill_2 FILLER_20_844 ();
 sg13g2_fill_1 FILLER_20_846 ();
 sg13g2_fill_1 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_20_883 ();
 sg13g2_decap_8 FILLER_20_890 ();
 sg13g2_fill_2 FILLER_20_897 ();
 sg13g2_fill_1 FILLER_20_899 ();
 sg13g2_decap_8 FILLER_20_914 ();
 sg13g2_decap_8 FILLER_20_921 ();
 sg13g2_decap_8 FILLER_20_928 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_decap_8 FILLER_20_942 ();
 sg13g2_decap_8 FILLER_20_949 ();
 sg13g2_decap_8 FILLER_20_956 ();
 sg13g2_decap_8 FILLER_20_963 ();
 sg13g2_decap_8 FILLER_20_970 ();
 sg13g2_decap_8 FILLER_20_977 ();
 sg13g2_decap_8 FILLER_20_984 ();
 sg13g2_decap_8 FILLER_20_991 ();
 sg13g2_decap_8 FILLER_20_998 ();
 sg13g2_decap_8 FILLER_20_1005 ();
 sg13g2_decap_8 FILLER_20_1012 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_decap_4 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_decap_4 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_93 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_4 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_decap_4 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_4 FILLER_21_378 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_1 FILLER_21_430 ();
 sg13g2_decap_8 FILLER_21_435 ();
 sg13g2_decap_8 FILLER_21_442 ();
 sg13g2_decap_8 FILLER_21_449 ();
 sg13g2_decap_4 FILLER_21_456 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_fill_2 FILLER_21_476 ();
 sg13g2_fill_1 FILLER_21_478 ();
 sg13g2_fill_1 FILLER_21_496 ();
 sg13g2_decap_8 FILLER_21_507 ();
 sg13g2_decap_4 FILLER_21_514 ();
 sg13g2_decap_4 FILLER_21_528 ();
 sg13g2_fill_1 FILLER_21_532 ();
 sg13g2_fill_1 FILLER_21_537 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_4 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_596 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_fill_1 FILLER_21_652 ();
 sg13g2_fill_2 FILLER_21_657 ();
 sg13g2_fill_2 FILLER_21_691 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_757 ();
 sg13g2_fill_2 FILLER_21_764 ();
 sg13g2_fill_1 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_4 FILLER_21_800 ();
 sg13g2_fill_1 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_813 ();
 sg13g2_decap_8 FILLER_21_820 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_fill_2 FILLER_21_849 ();
 sg13g2_decap_8 FILLER_21_870 ();
 sg13g2_decap_8 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_21_884 ();
 sg13g2_decap_8 FILLER_21_891 ();
 sg13g2_decap_4 FILLER_21_898 ();
 sg13g2_fill_1 FILLER_21_902 ();
 sg13g2_decap_8 FILLER_21_908 ();
 sg13g2_decap_8 FILLER_21_915 ();
 sg13g2_decap_8 FILLER_21_922 ();
 sg13g2_decap_8 FILLER_21_929 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_950 ();
 sg13g2_decap_8 FILLER_21_957 ();
 sg13g2_decap_8 FILLER_21_964 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_decap_8 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_985 ();
 sg13g2_decap_8 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_999 ();
 sg13g2_decap_8 FILLER_21_1006 ();
 sg13g2_decap_8 FILLER_21_1013 ();
 sg13g2_decap_8 FILLER_21_1020 ();
 sg13g2_fill_2 FILLER_21_1027 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_4 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_8 FILLER_22_78 ();
 sg13g2_decap_8 FILLER_22_85 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_decap_4 FILLER_22_417 ();
 sg13g2_fill_2 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_477 ();
 sg13g2_fill_2 FILLER_22_516 ();
 sg13g2_decap_8 FILLER_22_555 ();
 sg13g2_decap_8 FILLER_22_562 ();
 sg13g2_decap_8 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_576 ();
 sg13g2_decap_4 FILLER_22_583 ();
 sg13g2_decap_8 FILLER_22_619 ();
 sg13g2_decap_8 FILLER_22_626 ();
 sg13g2_decap_4 FILLER_22_633 ();
 sg13g2_decap_8 FILLER_22_645 ();
 sg13g2_fill_1 FILLER_22_652 ();
 sg13g2_decap_8 FILLER_22_675 ();
 sg13g2_fill_1 FILLER_22_682 ();
 sg13g2_fill_2 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_708 ();
 sg13g2_decap_8 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_722 ();
 sg13g2_decap_4 FILLER_22_729 ();
 sg13g2_fill_1 FILLER_22_733 ();
 sg13g2_decap_8 FILLER_22_754 ();
 sg13g2_decap_8 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_768 ();
 sg13g2_fill_2 FILLER_22_775 ();
 sg13g2_decap_8 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_789 ();
 sg13g2_decap_8 FILLER_22_796 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_decap_8 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_838 ();
 sg13g2_fill_1 FILLER_22_845 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_decap_8 FILLER_22_921 ();
 sg13g2_decap_8 FILLER_22_928 ();
 sg13g2_decap_8 FILLER_22_935 ();
 sg13g2_decap_8 FILLER_22_942 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_956 ();
 sg13g2_decap_8 FILLER_22_963 ();
 sg13g2_decap_8 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_decap_8 FILLER_22_991 ();
 sg13g2_decap_8 FILLER_22_998 ();
 sg13g2_decap_8 FILLER_22_1005 ();
 sg13g2_decap_8 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1019 ();
 sg13g2_fill_2 FILLER_22_1026 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_20 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_4 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_decap_4 FILLER_23_368 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_decap_4 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_435 ();
 sg13g2_decap_8 FILLER_23_442 ();
 sg13g2_fill_2 FILLER_23_449 ();
 sg13g2_decap_4 FILLER_23_455 ();
 sg13g2_fill_1 FILLER_23_459 ();
 sg13g2_fill_2 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_481 ();
 sg13g2_decap_4 FILLER_23_488 ();
 sg13g2_fill_2 FILLER_23_492 ();
 sg13g2_fill_2 FILLER_23_498 ();
 sg13g2_fill_1 FILLER_23_500 ();
 sg13g2_fill_2 FILLER_23_505 ();
 sg13g2_fill_2 FILLER_23_534 ();
 sg13g2_fill_1 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_541 ();
 sg13g2_decap_8 FILLER_23_548 ();
 sg13g2_decap_8 FILLER_23_555 ();
 sg13g2_decap_8 FILLER_23_562 ();
 sg13g2_decap_8 FILLER_23_569 ();
 sg13g2_fill_1 FILLER_23_576 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_597 ();
 sg13g2_decap_8 FILLER_23_604 ();
 sg13g2_decap_8 FILLER_23_611 ();
 sg13g2_decap_8 FILLER_23_618 ();
 sg13g2_decap_8 FILLER_23_625 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_4 FILLER_23_679 ();
 sg13g2_fill_1 FILLER_23_683 ();
 sg13g2_fill_2 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_727 ();
 sg13g2_fill_2 FILLER_23_734 ();
 sg13g2_fill_1 FILLER_23_736 ();
 sg13g2_decap_8 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_757 ();
 sg13g2_fill_1 FILLER_23_764 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_fill_2 FILLER_23_840 ();
 sg13g2_fill_1 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_871 ();
 sg13g2_decap_8 FILLER_23_878 ();
 sg13g2_decap_8 FILLER_23_885 ();
 sg13g2_decap_8 FILLER_23_892 ();
 sg13g2_decap_8 FILLER_23_899 ();
 sg13g2_decap_8 FILLER_23_906 ();
 sg13g2_decap_8 FILLER_23_913 ();
 sg13g2_decap_8 FILLER_23_920 ();
 sg13g2_decap_8 FILLER_23_927 ();
 sg13g2_decap_8 FILLER_23_934 ();
 sg13g2_decap_8 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_948 ();
 sg13g2_decap_8 FILLER_23_955 ();
 sg13g2_decap_8 FILLER_23_962 ();
 sg13g2_decap_8 FILLER_23_969 ();
 sg13g2_decap_8 FILLER_23_976 ();
 sg13g2_decap_8 FILLER_23_983 ();
 sg13g2_decap_8 FILLER_23_990 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_decap_8 FILLER_23_1004 ();
 sg13g2_decap_8 FILLER_23_1011 ();
 sg13g2_decap_8 FILLER_23_1018 ();
 sg13g2_decap_4 FILLER_23_1025 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_38 ();
 sg13g2_decap_4 FILLER_24_45 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_4 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_fill_1 FILLER_24_400 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_fill_1 FILLER_24_425 ();
 sg13g2_decap_4 FILLER_24_453 ();
 sg13g2_fill_1 FILLER_24_457 ();
 sg13g2_decap_4 FILLER_24_466 ();
 sg13g2_fill_1 FILLER_24_470 ();
 sg13g2_decap_8 FILLER_24_485 ();
 sg13g2_decap_8 FILLER_24_506 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_4 FILLER_24_567 ();
 sg13g2_fill_1 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_decap_4 FILLER_24_642 ();
 sg13g2_fill_1 FILLER_24_646 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_fill_2 FILLER_24_681 ();
 sg13g2_fill_1 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_fill_2 FILLER_24_754 ();
 sg13g2_fill_1 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_fill_2 FILLER_24_791 ();
 sg13g2_fill_1 FILLER_24_793 ();
 sg13g2_decap_4 FILLER_24_803 ();
 sg13g2_fill_1 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_4 FILLER_24_849 ();
 sg13g2_decap_8 FILLER_24_862 ();
 sg13g2_decap_8 FILLER_24_869 ();
 sg13g2_decap_8 FILLER_24_876 ();
 sg13g2_decap_8 FILLER_24_883 ();
 sg13g2_decap_8 FILLER_24_890 ();
 sg13g2_decap_8 FILLER_24_897 ();
 sg13g2_decap_8 FILLER_24_904 ();
 sg13g2_decap_8 FILLER_24_911 ();
 sg13g2_decap_8 FILLER_24_918 ();
 sg13g2_decap_8 FILLER_24_925 ();
 sg13g2_decap_8 FILLER_24_932 ();
 sg13g2_decap_8 FILLER_24_939 ();
 sg13g2_decap_8 FILLER_24_946 ();
 sg13g2_decap_8 FILLER_24_953 ();
 sg13g2_decap_8 FILLER_24_960 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_decap_8 FILLER_24_981 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_decap_8 FILLER_24_995 ();
 sg13g2_decap_8 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1009 ();
 sg13g2_decap_8 FILLER_24_1016 ();
 sg13g2_decap_4 FILLER_24_1023 ();
 sg13g2_fill_2 FILLER_24_1027 ();
 sg13g2_fill_2 FILLER_25_20 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_decap_4 FILLER_25_51 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_4 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_4 FILLER_25_358 ();
 sg13g2_decap_4 FILLER_25_393 ();
 sg13g2_decap_4 FILLER_25_401 ();
 sg13g2_fill_2 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_420 ();
 sg13g2_decap_4 FILLER_25_447 ();
 sg13g2_fill_2 FILLER_25_451 ();
 sg13g2_fill_2 FILLER_25_484 ();
 sg13g2_fill_1 FILLER_25_492 ();
 sg13g2_decap_4 FILLER_25_507 ();
 sg13g2_fill_1 FILLER_25_511 ();
 sg13g2_decap_4 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_535 ();
 sg13g2_fill_2 FILLER_25_542 ();
 sg13g2_decap_4 FILLER_25_549 ();
 sg13g2_fill_1 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_decap_4 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_593 ();
 sg13g2_decap_8 FILLER_25_598 ();
 sg13g2_decap_4 FILLER_25_605 ();
 sg13g2_fill_2 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_628 ();
 sg13g2_decap_8 FILLER_25_635 ();
 sg13g2_decap_8 FILLER_25_642 ();
 sg13g2_fill_2 FILLER_25_649 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_fill_2 FILLER_25_748 ();
 sg13g2_fill_1 FILLER_25_750 ();
 sg13g2_decap_4 FILLER_25_781 ();
 sg13g2_fill_1 FILLER_25_785 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_2 FILLER_25_807 ();
 sg13g2_fill_1 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_fill_1 FILLER_25_830 ();
 sg13g2_decap_4 FILLER_25_836 ();
 sg13g2_fill_2 FILLER_25_847 ();
 sg13g2_fill_1 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_871 ();
 sg13g2_decap_8 FILLER_25_878 ();
 sg13g2_decap_8 FILLER_25_885 ();
 sg13g2_decap_8 FILLER_25_892 ();
 sg13g2_decap_8 FILLER_25_899 ();
 sg13g2_decap_8 FILLER_25_906 ();
 sg13g2_decap_8 FILLER_25_913 ();
 sg13g2_decap_8 FILLER_25_920 ();
 sg13g2_decap_8 FILLER_25_927 ();
 sg13g2_decap_8 FILLER_25_934 ();
 sg13g2_decap_8 FILLER_25_941 ();
 sg13g2_decap_8 FILLER_25_948 ();
 sg13g2_decap_8 FILLER_25_955 ();
 sg13g2_decap_8 FILLER_25_962 ();
 sg13g2_decap_8 FILLER_25_969 ();
 sg13g2_decap_8 FILLER_25_976 ();
 sg13g2_decap_8 FILLER_25_983 ();
 sg13g2_decap_8 FILLER_25_990 ();
 sg13g2_decap_8 FILLER_25_997 ();
 sg13g2_decap_8 FILLER_25_1004 ();
 sg13g2_decap_8 FILLER_25_1011 ();
 sg13g2_decap_8 FILLER_25_1018 ();
 sg13g2_decap_4 FILLER_25_1025 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_decap_4 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_44 ();
 sg13g2_decap_4 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_55 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_75 ();
 sg13g2_decap_8 FILLER_26_82 ();
 sg13g2_decap_4 FILLER_26_89 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_4 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_284 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_decap_4 FILLER_26_392 ();
 sg13g2_fill_2 FILLER_26_433 ();
 sg13g2_fill_1 FILLER_26_435 ();
 sg13g2_decap_4 FILLER_26_449 ();
 sg13g2_fill_2 FILLER_26_470 ();
 sg13g2_fill_1 FILLER_26_472 ();
 sg13g2_decap_8 FILLER_26_478 ();
 sg13g2_decap_8 FILLER_26_485 ();
 sg13g2_fill_1 FILLER_26_492 ();
 sg13g2_decap_8 FILLER_26_510 ();
 sg13g2_decap_8 FILLER_26_522 ();
 sg13g2_decap_8 FILLER_26_529 ();
 sg13g2_fill_2 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_575 ();
 sg13g2_decap_8 FILLER_26_582 ();
 sg13g2_decap_8 FILLER_26_629 ();
 sg13g2_decap_8 FILLER_26_636 ();
 sg13g2_decap_8 FILLER_26_643 ();
 sg13g2_fill_2 FILLER_26_650 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_fill_1 FILLER_26_684 ();
 sg13g2_fill_2 FILLER_26_694 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_1 FILLER_26_738 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_4 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_766 ();
 sg13g2_decap_4 FILLER_26_773 ();
 sg13g2_fill_2 FILLER_26_777 ();
 sg13g2_fill_1 FILLER_26_792 ();
 sg13g2_fill_1 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_fill_2 FILLER_26_822 ();
 sg13g2_fill_1 FILLER_26_824 ();
 sg13g2_fill_1 FILLER_26_857 ();
 sg13g2_fill_2 FILLER_26_868 ();
 sg13g2_fill_1 FILLER_26_870 ();
 sg13g2_decap_8 FILLER_26_884 ();
 sg13g2_decap_8 FILLER_26_891 ();
 sg13g2_decap_8 FILLER_26_898 ();
 sg13g2_decap_8 FILLER_26_905 ();
 sg13g2_decap_8 FILLER_26_912 ();
 sg13g2_decap_8 FILLER_26_919 ();
 sg13g2_decap_8 FILLER_26_926 ();
 sg13g2_decap_8 FILLER_26_933 ();
 sg13g2_decap_8 FILLER_26_940 ();
 sg13g2_decap_8 FILLER_26_947 ();
 sg13g2_decap_8 FILLER_26_954 ();
 sg13g2_decap_8 FILLER_26_961 ();
 sg13g2_decap_8 FILLER_26_968 ();
 sg13g2_decap_8 FILLER_26_975 ();
 sg13g2_decap_8 FILLER_26_982 ();
 sg13g2_decap_8 FILLER_26_989 ();
 sg13g2_decap_8 FILLER_26_996 ();
 sg13g2_decap_8 FILLER_26_1003 ();
 sg13g2_decap_8 FILLER_26_1010 ();
 sg13g2_decap_8 FILLER_26_1017 ();
 sg13g2_decap_4 FILLER_26_1024 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_6 ();
 sg13g2_decap_4 FILLER_27_11 ();
 sg13g2_decap_8 FILLER_27_19 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_fill_2 FILLER_27_48 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_decap_4 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_decap_4 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_410 ();
 sg13g2_fill_1 FILLER_27_412 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_4 FILLER_27_435 ();
 sg13g2_fill_1 FILLER_27_439 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_464 ();
 sg13g2_fill_1 FILLER_27_486 ();
 sg13g2_fill_2 FILLER_27_537 ();
 sg13g2_decap_4 FILLER_27_542 ();
 sg13g2_fill_2 FILLER_27_546 ();
 sg13g2_fill_2 FILLER_27_552 ();
 sg13g2_fill_2 FILLER_27_558 ();
 sg13g2_decap_8 FILLER_27_565 ();
 sg13g2_decap_8 FILLER_27_572 ();
 sg13g2_decap_8 FILLER_27_579 ();
 sg13g2_decap_8 FILLER_27_586 ();
 sg13g2_decap_8 FILLER_27_593 ();
 sg13g2_decap_8 FILLER_27_600 ();
 sg13g2_decap_4 FILLER_27_607 ();
 sg13g2_decap_8 FILLER_27_615 ();
 sg13g2_fill_2 FILLER_27_622 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_decap_4 FILLER_27_638 ();
 sg13g2_fill_2 FILLER_27_654 ();
 sg13g2_decap_4 FILLER_27_661 ();
 sg13g2_decap_4 FILLER_27_675 ();
 sg13g2_fill_1 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_708 ();
 sg13g2_decap_8 FILLER_27_715 ();
 sg13g2_decap_4 FILLER_27_722 ();
 sg13g2_fill_2 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_fill_2 FILLER_27_786 ();
 sg13g2_fill_1 FILLER_27_788 ();
 sg13g2_decap_8 FILLER_27_806 ();
 sg13g2_decap_4 FILLER_27_813 ();
 sg13g2_fill_2 FILLER_27_826 ();
 sg13g2_fill_1 FILLER_27_828 ();
 sg13g2_decap_4 FILLER_27_850 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_29 ();
 sg13g2_decap_8 FILLER_28_36 ();
 sg13g2_decap_8 FILLER_28_43 ();
 sg13g2_decap_4 FILLER_28_50 ();
 sg13g2_decap_4 FILLER_28_68 ();
 sg13g2_decap_8 FILLER_28_93 ();
 sg13g2_decap_8 FILLER_28_100 ();
 sg13g2_fill_2 FILLER_28_107 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_decap_4 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_decap_4 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_431 ();
 sg13g2_decap_8 FILLER_28_446 ();
 sg13g2_decap_8 FILLER_28_453 ();
 sg13g2_fill_1 FILLER_28_460 ();
 sg13g2_decap_8 FILLER_28_474 ();
 sg13g2_decap_8 FILLER_28_481 ();
 sg13g2_decap_8 FILLER_28_488 ();
 sg13g2_fill_2 FILLER_28_495 ();
 sg13g2_fill_1 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_502 ();
 sg13g2_decap_8 FILLER_28_509 ();
 sg13g2_fill_2 FILLER_28_516 ();
 sg13g2_fill_1 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_fill_1 FILLER_28_531 ();
 sg13g2_fill_2 FILLER_28_550 ();
 sg13g2_fill_1 FILLER_28_552 ();
 sg13g2_fill_2 FILLER_28_560 ();
 sg13g2_fill_1 FILLER_28_562 ();
 sg13g2_decap_8 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_597 ();
 sg13g2_fill_2 FILLER_28_604 ();
 sg13g2_decap_4 FILLER_28_633 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_fill_2 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_4 FILLER_28_699 ();
 sg13g2_fill_2 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_709 ();
 sg13g2_decap_8 FILLER_28_716 ();
 sg13g2_decap_4 FILLER_28_723 ();
 sg13g2_fill_1 FILLER_28_727 ();
 sg13g2_fill_1 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_fill_1 FILLER_28_755 ();
 sg13g2_decap_4 FILLER_28_769 ();
 sg13g2_fill_1 FILLER_28_773 ();
 sg13g2_fill_1 FILLER_28_790 ();
 sg13g2_decap_4 FILLER_28_804 ();
 sg13g2_fill_2 FILLER_28_808 ();
 sg13g2_fill_1 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_fill_2 FILLER_28_852 ();
 sg13g2_fill_1 FILLER_28_854 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_8 FILLER_28_886 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_decap_8 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_935 ();
 sg13g2_decap_8 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_956 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_fill_2 FILLER_28_1026 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_fill_2 FILLER_29_5 ();
 sg13g2_decap_4 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_19 ();
 sg13g2_decap_8 FILLER_29_31 ();
 sg13g2_fill_2 FILLER_29_38 ();
 sg13g2_decap_8 FILLER_29_57 ();
 sg13g2_decap_8 FILLER_29_64 ();
 sg13g2_decap_8 FILLER_29_71 ();
 sg13g2_decap_8 FILLER_29_78 ();
 sg13g2_decap_8 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_29_409 ();
 sg13g2_fill_2 FILLER_29_416 ();
 sg13g2_fill_1 FILLER_29_418 ();
 sg13g2_decap_4 FILLER_29_459 ();
 sg13g2_fill_1 FILLER_29_463 ();
 sg13g2_fill_2 FILLER_29_491 ();
 sg13g2_fill_2 FILLER_29_509 ();
 sg13g2_decap_8 FILLER_29_538 ();
 sg13g2_decap_4 FILLER_29_555 ();
 sg13g2_decap_4 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_572 ();
 sg13g2_decap_8 FILLER_29_579 ();
 sg13g2_decap_8 FILLER_29_586 ();
 sg13g2_decap_8 FILLER_29_593 ();
 sg13g2_decap_4 FILLER_29_600 ();
 sg13g2_fill_2 FILLER_29_604 ();
 sg13g2_fill_1 FILLER_29_611 ();
 sg13g2_decap_8 FILLER_29_617 ();
 sg13g2_fill_2 FILLER_29_624 ();
 sg13g2_fill_2 FILLER_29_645 ();
 sg13g2_fill_2 FILLER_29_656 ();
 sg13g2_fill_1 FILLER_29_658 ();
 sg13g2_fill_2 FILLER_29_663 ();
 sg13g2_fill_1 FILLER_29_665 ();
 sg13g2_decap_4 FILLER_29_675 ();
 sg13g2_decap_4 FILLER_29_724 ();
 sg13g2_fill_1 FILLER_29_728 ();
 sg13g2_decap_4 FILLER_29_737 ();
 sg13g2_fill_1 FILLER_29_741 ();
 sg13g2_fill_2 FILLER_29_750 ();
 sg13g2_fill_1 FILLER_29_752 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_4 FILLER_29_772 ();
 sg13g2_fill_1 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_796 ();
 sg13g2_decap_8 FILLER_29_803 ();
 sg13g2_decap_4 FILLER_29_810 ();
 sg13g2_fill_2 FILLER_29_848 ();
 sg13g2_fill_1 FILLER_29_850 ();
 sg13g2_fill_2 FILLER_29_855 ();
 sg13g2_decap_8 FILLER_29_890 ();
 sg13g2_decap_8 FILLER_29_897 ();
 sg13g2_decap_8 FILLER_29_904 ();
 sg13g2_decap_8 FILLER_29_911 ();
 sg13g2_decap_8 FILLER_29_918 ();
 sg13g2_decap_8 FILLER_29_925 ();
 sg13g2_decap_8 FILLER_29_932 ();
 sg13g2_decap_8 FILLER_29_939 ();
 sg13g2_decap_8 FILLER_29_946 ();
 sg13g2_decap_8 FILLER_29_953 ();
 sg13g2_decap_8 FILLER_29_960 ();
 sg13g2_decap_8 FILLER_29_967 ();
 sg13g2_decap_8 FILLER_29_974 ();
 sg13g2_decap_8 FILLER_29_981 ();
 sg13g2_decap_8 FILLER_29_988 ();
 sg13g2_decap_8 FILLER_29_995 ();
 sg13g2_decap_8 FILLER_29_1002 ();
 sg13g2_decap_8 FILLER_29_1009 ();
 sg13g2_decap_8 FILLER_29_1016 ();
 sg13g2_decap_4 FILLER_29_1023 ();
 sg13g2_fill_2 FILLER_29_1027 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_decap_4 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_decap_4 FILLER_30_395 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_417 ();
 sg13g2_fill_1 FILLER_30_419 ();
 sg13g2_fill_1 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_439 ();
 sg13g2_fill_1 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_447 ();
 sg13g2_decap_4 FILLER_30_454 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_decap_4 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_481 ();
 sg13g2_decap_4 FILLER_30_496 ();
 sg13g2_fill_1 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_505 ();
 sg13g2_fill_2 FILLER_30_520 ();
 sg13g2_decap_8 FILLER_30_526 ();
 sg13g2_decap_8 FILLER_30_533 ();
 sg13g2_decap_4 FILLER_30_540 ();
 sg13g2_fill_2 FILLER_30_544 ();
 sg13g2_decap_8 FILLER_30_578 ();
 sg13g2_decap_8 FILLER_30_585 ();
 sg13g2_fill_1 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_2 FILLER_30_620 ();
 sg13g2_fill_2 FILLER_30_640 ();
 sg13g2_fill_1 FILLER_30_642 ();
 sg13g2_fill_2 FILLER_30_663 ();
 sg13g2_decap_4 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_703 ();
 sg13g2_decap_8 FILLER_30_710 ();
 sg13g2_fill_2 FILLER_30_717 ();
 sg13g2_fill_1 FILLER_30_719 ();
 sg13g2_fill_1 FILLER_30_747 ();
 sg13g2_decap_4 FILLER_30_769 ();
 sg13g2_fill_2 FILLER_30_787 ();
 sg13g2_fill_2 FILLER_30_821 ();
 sg13g2_fill_2 FILLER_30_827 ();
 sg13g2_fill_1 FILLER_30_829 ();
 sg13g2_decap_8 FILLER_30_845 ();
 sg13g2_decap_8 FILLER_30_852 ();
 sg13g2_decap_4 FILLER_30_859 ();
 sg13g2_fill_2 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_874 ();
 sg13g2_decap_8 FILLER_30_881 ();
 sg13g2_decap_8 FILLER_30_888 ();
 sg13g2_decap_8 FILLER_30_895 ();
 sg13g2_decap_8 FILLER_30_902 ();
 sg13g2_decap_8 FILLER_30_909 ();
 sg13g2_decap_8 FILLER_30_916 ();
 sg13g2_decap_8 FILLER_30_923 ();
 sg13g2_decap_8 FILLER_30_930 ();
 sg13g2_decap_8 FILLER_30_937 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_decap_8 FILLER_30_951 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_decap_8 FILLER_30_965 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_986 ();
 sg13g2_decap_8 FILLER_30_993 ();
 sg13g2_decap_8 FILLER_30_1000 ();
 sg13g2_decap_8 FILLER_30_1007 ();
 sg13g2_decap_8 FILLER_30_1014 ();
 sg13g2_decap_8 FILLER_30_1021 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_8 FILLER_31_5 ();
 sg13g2_decap_8 FILLER_31_12 ();
 sg13g2_fill_2 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_4 FILLER_31_395 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_428 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_fill_2 FILLER_31_441 ();
 sg13g2_fill_1 FILLER_31_443 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_459 ();
 sg13g2_fill_2 FILLER_31_466 ();
 sg13g2_fill_2 FILLER_31_481 ();
 sg13g2_fill_2 FILLER_31_510 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_fill_2 FILLER_31_581 ();
 sg13g2_fill_1 FILLER_31_583 ();
 sg13g2_decap_8 FILLER_31_614 ();
 sg13g2_decap_8 FILLER_31_621 ();
 sg13g2_decap_4 FILLER_31_640 ();
 sg13g2_fill_2 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_fill_2 FILLER_31_693 ();
 sg13g2_fill_1 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_723 ();
 sg13g2_decap_8 FILLER_31_747 ();
 sg13g2_fill_1 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_fill_1 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_837 ();
 sg13g2_decap_8 FILLER_31_899 ();
 sg13g2_decap_8 FILLER_31_906 ();
 sg13g2_decap_8 FILLER_31_913 ();
 sg13g2_decap_8 FILLER_31_920 ();
 sg13g2_decap_8 FILLER_31_927 ();
 sg13g2_decap_8 FILLER_31_934 ();
 sg13g2_decap_8 FILLER_31_941 ();
 sg13g2_decap_8 FILLER_31_948 ();
 sg13g2_decap_8 FILLER_31_955 ();
 sg13g2_decap_8 FILLER_31_962 ();
 sg13g2_decap_8 FILLER_31_969 ();
 sg13g2_decap_8 FILLER_31_976 ();
 sg13g2_decap_8 FILLER_31_983 ();
 sg13g2_decap_8 FILLER_31_990 ();
 sg13g2_decap_8 FILLER_31_997 ();
 sg13g2_decap_8 FILLER_31_1004 ();
 sg13g2_decap_8 FILLER_31_1011 ();
 sg13g2_decap_8 FILLER_31_1018 ();
 sg13g2_decap_4 FILLER_31_1025 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_40 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_decap_4 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_decap_4 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_decap_4 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_4 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_366 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_decap_4 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_fill_1 FILLER_32_417 ();
 sg13g2_fill_1 FILLER_32_423 ();
 sg13g2_decap_4 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_510 ();
 sg13g2_decap_8 FILLER_32_521 ();
 sg13g2_decap_8 FILLER_32_528 ();
 sg13g2_decap_4 FILLER_32_535 ();
 sg13g2_fill_2 FILLER_32_539 ();
 sg13g2_fill_1 FILLER_32_548 ();
 sg13g2_decap_8 FILLER_32_576 ();
 sg13g2_decap_8 FILLER_32_583 ();
 sg13g2_fill_2 FILLER_32_590 ();
 sg13g2_fill_2 FILLER_32_596 ();
 sg13g2_decap_8 FILLER_32_625 ();
 sg13g2_decap_8 FILLER_32_632 ();
 sg13g2_decap_8 FILLER_32_639 ();
 sg13g2_decap_4 FILLER_32_646 ();
 sg13g2_fill_2 FILLER_32_654 ();
 sg13g2_fill_1 FILLER_32_656 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_decap_4 FILLER_32_675 ();
 sg13g2_fill_2 FILLER_32_679 ();
 sg13g2_fill_2 FILLER_32_689 ();
 sg13g2_fill_1 FILLER_32_691 ();
 sg13g2_fill_1 FILLER_32_698 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_8 FILLER_32_715 ();
 sg13g2_fill_1 FILLER_32_737 ();
 sg13g2_decap_8 FILLER_32_765 ();
 sg13g2_decap_8 FILLER_32_772 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_4 FILLER_32_824 ();
 sg13g2_decap_8 FILLER_32_860 ();
 sg13g2_decap_4 FILLER_32_867 ();
 sg13g2_decap_8 FILLER_32_902 ();
 sg13g2_decap_8 FILLER_32_909 ();
 sg13g2_decap_8 FILLER_32_916 ();
 sg13g2_decap_8 FILLER_32_923 ();
 sg13g2_decap_8 FILLER_32_930 ();
 sg13g2_decap_8 FILLER_32_937 ();
 sg13g2_decap_8 FILLER_32_948 ();
 sg13g2_decap_8 FILLER_32_955 ();
 sg13g2_decap_8 FILLER_32_962 ();
 sg13g2_decap_8 FILLER_32_969 ();
 sg13g2_decap_8 FILLER_32_976 ();
 sg13g2_decap_8 FILLER_32_983 ();
 sg13g2_decap_8 FILLER_32_990 ();
 sg13g2_decap_8 FILLER_32_997 ();
 sg13g2_decap_8 FILLER_32_1004 ();
 sg13g2_decap_8 FILLER_32_1011 ();
 sg13g2_decap_8 FILLER_32_1018 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_1 FILLER_33_13 ();
 sg13g2_decap_4 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_22 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_decap_4 FILLER_33_72 ();
 sg13g2_fill_2 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_decap_4 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_4 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_decap_4 FILLER_33_430 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_439 ();
 sg13g2_fill_2 FILLER_33_445 ();
 sg13g2_decap_4 FILLER_33_451 ();
 sg13g2_decap_4 FILLER_33_465 ();
 sg13g2_fill_2 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_475 ();
 sg13g2_decap_4 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_486 ();
 sg13g2_decap_4 FILLER_33_492 ();
 sg13g2_fill_1 FILLER_33_496 ();
 sg13g2_decap_4 FILLER_33_510 ();
 sg13g2_fill_1 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_519 ();
 sg13g2_decap_8 FILLER_33_526 ();
 sg13g2_fill_2 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_607 ();
 sg13g2_decap_4 FILLER_33_614 ();
 sg13g2_fill_1 FILLER_33_618 ();
 sg13g2_fill_2 FILLER_33_734 ();
 sg13g2_decap_4 FILLER_33_782 ();
 sg13g2_fill_2 FILLER_33_786 ();
 sg13g2_decap_4 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_4 FILLER_33_813 ();
 sg13g2_fill_1 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_4 FILLER_33_859 ();
 sg13g2_fill_2 FILLER_33_863 ();
 sg13g2_fill_2 FILLER_33_878 ();
 sg13g2_decap_8 FILLER_33_884 ();
 sg13g2_decap_4 FILLER_33_891 ();
 sg13g2_fill_1 FILLER_33_895 ();
 sg13g2_decap_8 FILLER_33_901 ();
 sg13g2_fill_2 FILLER_33_908 ();
 sg13g2_fill_1 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_4 FILLER_33_931 ();
 sg13g2_fill_2 FILLER_33_947 ();
 sg13g2_decap_8 FILLER_33_958 ();
 sg13g2_decap_8 FILLER_33_965 ();
 sg13g2_decap_8 FILLER_33_972 ();
 sg13g2_decap_8 FILLER_33_979 ();
 sg13g2_decap_8 FILLER_33_986 ();
 sg13g2_decap_8 FILLER_33_993 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_decap_8 FILLER_33_1007 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_decap_4 FILLER_34_9 ();
 sg13g2_fill_1 FILLER_34_17 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_decap_8 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_decap_8 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_decap_4 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_325 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_decap_4 FILLER_34_349 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_419 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_fill_1 FILLER_34_459 ();
 sg13g2_decap_4 FILLER_34_487 ();
 sg13g2_fill_1 FILLER_34_501 ();
 sg13g2_decap_8 FILLER_34_529 ();
 sg13g2_decap_4 FILLER_34_536 ();
 sg13g2_decap_4 FILLER_34_544 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_568 ();
 sg13g2_decap_8 FILLER_34_578 ();
 sg13g2_fill_2 FILLER_34_585 ();
 sg13g2_decap_4 FILLER_34_619 ();
 sg13g2_fill_1 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_fill_2 FILLER_34_651 ();
 sg13g2_fill_1 FILLER_34_653 ();
 sg13g2_fill_2 FILLER_34_682 ();
 sg13g2_fill_1 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_689 ();
 sg13g2_decap_8 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_703 ();
 sg13g2_decap_8 FILLER_34_710 ();
 sg13g2_decap_8 FILLER_34_717 ();
 sg13g2_decap_8 FILLER_34_724 ();
 sg13g2_fill_1 FILLER_34_731 ();
 sg13g2_decap_8 FILLER_34_745 ();
 sg13g2_decap_4 FILLER_34_752 ();
 sg13g2_decap_4 FILLER_34_764 ();
 sg13g2_fill_2 FILLER_34_795 ();
 sg13g2_fill_1 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_844 ();
 sg13g2_decap_8 FILLER_34_851 ();
 sg13g2_decap_8 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_34_865 ();
 sg13g2_fill_2 FILLER_34_872 ();
 sg13g2_decap_8 FILLER_34_879 ();
 sg13g2_decap_4 FILLER_34_886 ();
 sg13g2_fill_2 FILLER_34_898 ();
 sg13g2_decap_8 FILLER_34_921 ();
 sg13g2_fill_1 FILLER_34_928 ();
 sg13g2_fill_1 FILLER_34_945 ();
 sg13g2_fill_2 FILLER_34_954 ();
 sg13g2_fill_1 FILLER_34_956 ();
 sg13g2_decap_8 FILLER_34_972 ();
 sg13g2_decap_8 FILLER_34_979 ();
 sg13g2_decap_8 FILLER_34_986 ();
 sg13g2_decap_8 FILLER_34_993 ();
 sg13g2_decap_8 FILLER_34_1000 ();
 sg13g2_decap_8 FILLER_34_1007 ();
 sg13g2_decap_8 FILLER_34_1014 ();
 sg13g2_decap_8 FILLER_34_1021 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_72 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_decap_8 FILLER_35_121 ();
 sg13g2_fill_2 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_decap_4 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_decap_4 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_decap_4 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_decap_4 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_decap_4 FILLER_35_390 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_438 ();
 sg13g2_decap_8 FILLER_35_445 ();
 sg13g2_fill_1 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_463 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_4 FILLER_35_483 ();
 sg13g2_fill_2 FILLER_35_487 ();
 sg13g2_fill_2 FILLER_35_506 ();
 sg13g2_fill_2 FILLER_35_512 ();
 sg13g2_fill_1 FILLER_35_514 ();
 sg13g2_fill_2 FILLER_35_519 ();
 sg13g2_fill_1 FILLER_35_521 ();
 sg13g2_decap_8 FILLER_35_526 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_fill_1 FILLER_35_540 ();
 sg13g2_decap_4 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_577 ();
 sg13g2_fill_1 FILLER_35_579 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_fill_1 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_599 ();
 sg13g2_decap_4 FILLER_35_606 ();
 sg13g2_fill_2 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_628 ();
 sg13g2_decap_4 FILLER_35_633 ();
 sg13g2_fill_1 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_642 ();
 sg13g2_decap_8 FILLER_35_649 ();
 sg13g2_fill_2 FILLER_35_656 ();
 sg13g2_fill_1 FILLER_35_658 ();
 sg13g2_fill_1 FILLER_35_663 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_8 FILLER_35_675 ();
 sg13g2_fill_1 FILLER_35_682 ();
 sg13g2_decap_4 FILLER_35_710 ();
 sg13g2_fill_2 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_fill_1 FILLER_35_757 ();
 sg13g2_decap_4 FILLER_35_766 ();
 sg13g2_fill_2 FILLER_35_770 ();
 sg13g2_decap_4 FILLER_35_817 ();
 sg13g2_fill_2 FILLER_35_821 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_4 FILLER_35_879 ();
 sg13g2_fill_2 FILLER_35_883 ();
 sg13g2_decap_4 FILLER_35_895 ();
 sg13g2_fill_2 FILLER_35_921 ();
 sg13g2_fill_2 FILLER_35_928 ();
 sg13g2_fill_1 FILLER_35_930 ();
 sg13g2_fill_1 FILLER_35_956 ();
 sg13g2_fill_1 FILLER_35_961 ();
 sg13g2_fill_2 FILLER_35_970 ();
 sg13g2_decap_8 FILLER_35_984 ();
 sg13g2_decap_8 FILLER_35_991 ();
 sg13g2_decap_8 FILLER_35_998 ();
 sg13g2_decap_8 FILLER_35_1005 ();
 sg13g2_decap_8 FILLER_35_1012 ();
 sg13g2_decap_8 FILLER_35_1019 ();
 sg13g2_fill_2 FILLER_35_1026 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_8 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_fill_2 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_decap_4 FILLER_36_414 ();
 sg13g2_fill_2 FILLER_36_418 ();
 sg13g2_fill_2 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_444 ();
 sg13g2_decap_4 FILLER_36_451 ();
 sg13g2_fill_1 FILLER_36_460 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_fill_2 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_537 ();
 sg13g2_decap_8 FILLER_36_544 ();
 sg13g2_decap_4 FILLER_36_551 ();
 sg13g2_fill_2 FILLER_36_555 ();
 sg13g2_fill_1 FILLER_36_578 ();
 sg13g2_fill_1 FILLER_36_584 ();
 sg13g2_decap_4 FILLER_36_590 ();
 sg13g2_fill_2 FILLER_36_594 ();
 sg13g2_decap_4 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_642 ();
 sg13g2_decap_4 FILLER_36_653 ();
 sg13g2_fill_2 FILLER_36_657 ();
 sg13g2_fill_2 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_698 ();
 sg13g2_fill_2 FILLER_36_705 ();
 sg13g2_fill_1 FILLER_36_707 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_fill_2 FILLER_36_868 ();
 sg13g2_fill_1 FILLER_36_870 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_fill_2 FILLER_36_886 ();
 sg13g2_decap_4 FILLER_36_894 ();
 sg13g2_decap_8 FILLER_36_921 ();
 sg13g2_fill_1 FILLER_36_928 ();
 sg13g2_fill_2 FILLER_36_938 ();
 sg13g2_fill_1 FILLER_36_940 ();
 sg13g2_decap_8 FILLER_36_946 ();
 sg13g2_decap_4 FILLER_36_953 ();
 sg13g2_fill_2 FILLER_36_957 ();
 sg13g2_fill_1 FILLER_36_970 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_50 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_fill_1 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_decap_4 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_decap_4 FILLER_37_157 ();
 sg13g2_decap_4 FILLER_37_192 ();
 sg13g2_decap_4 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_4 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_decap_4 FILLER_37_394 ();
 sg13g2_fill_1 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_412 ();
 sg13g2_fill_1 FILLER_37_447 ();
 sg13g2_decap_4 FILLER_37_489 ();
 sg13g2_fill_2 FILLER_37_512 ();
 sg13g2_fill_2 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_decap_8 FILLER_37_531 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_4 FILLER_37_545 ();
 sg13g2_fill_2 FILLER_37_568 ();
 sg13g2_fill_1 FILLER_37_570 ();
 sg13g2_fill_2 FILLER_37_584 ();
 sg13g2_fill_1 FILLER_37_586 ();
 sg13g2_decap_4 FILLER_37_593 ();
 sg13g2_fill_2 FILLER_37_597 ();
 sg13g2_fill_2 FILLER_37_604 ();
 sg13g2_decap_8 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_618 ();
 sg13g2_fill_1 FILLER_37_635 ();
 sg13g2_decap_8 FILLER_37_653 ();
 sg13g2_decap_8 FILLER_37_660 ();
 sg13g2_decap_8 FILLER_37_667 ();
 sg13g2_decap_8 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_fill_2 FILLER_37_720 ();
 sg13g2_decap_8 FILLER_37_726 ();
 sg13g2_decap_4 FILLER_37_733 ();
 sg13g2_fill_1 FILLER_37_737 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_fill_1 FILLER_37_755 ();
 sg13g2_fill_2 FILLER_37_810 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_4 FILLER_37_828 ();
 sg13g2_fill_2 FILLER_37_832 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_2 FILLER_37_876 ();
 sg13g2_fill_1 FILLER_37_878 ();
 sg13g2_decap_8 FILLER_37_884 ();
 sg13g2_decap_4 FILLER_37_891 ();
 sg13g2_decap_4 FILLER_37_921 ();
 sg13g2_fill_2 FILLER_37_951 ();
 sg13g2_fill_1 FILLER_37_953 ();
 sg13g2_decap_8 FILLER_37_983 ();
 sg13g2_decap_8 FILLER_37_990 ();
 sg13g2_decap_8 FILLER_37_997 ();
 sg13g2_decap_8 FILLER_37_1004 ();
 sg13g2_decap_8 FILLER_37_1011 ();
 sg13g2_decap_8 FILLER_37_1018 ();
 sg13g2_decap_4 FILLER_37_1025 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_53 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_4 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_fill_2 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_38_415 ();
 sg13g2_fill_2 FILLER_38_464 ();
 sg13g2_fill_1 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_471 ();
 sg13g2_decap_8 FILLER_38_478 ();
 sg13g2_decap_8 FILLER_38_500 ();
 sg13g2_fill_2 FILLER_38_507 ();
 sg13g2_decap_4 FILLER_38_536 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_decap_4 FILLER_38_574 ();
 sg13g2_fill_2 FILLER_38_578 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_decap_8 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_608 ();
 sg13g2_decap_8 FILLER_38_615 ();
 sg13g2_decap_4 FILLER_38_622 ();
 sg13g2_decap_4 FILLER_38_678 ();
 sg13g2_fill_2 FILLER_38_709 ();
 sg13g2_fill_1 FILLER_38_711 ();
 sg13g2_decap_4 FILLER_38_717 ();
 sg13g2_fill_2 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_4 FILLER_38_765 ();
 sg13g2_fill_2 FILLER_38_769 ();
 sg13g2_decap_4 FILLER_38_784 ();
 sg13g2_fill_1 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_4 FILLER_38_812 ();
 sg13g2_fill_2 FILLER_38_829 ();
 sg13g2_fill_1 FILLER_38_831 ();
 sg13g2_fill_2 FILLER_38_856 ();
 sg13g2_fill_1 FILLER_38_858 ();
 sg13g2_decap_4 FILLER_38_878 ();
 sg13g2_decap_4 FILLER_38_895 ();
 sg13g2_decap_8 FILLER_38_912 ();
 sg13g2_decap_8 FILLER_38_919 ();
 sg13g2_fill_1 FILLER_38_926 ();
 sg13g2_decap_8 FILLER_38_950 ();
 sg13g2_fill_2 FILLER_38_957 ();
 sg13g2_decap_8 FILLER_38_972 ();
 sg13g2_decap_8 FILLER_38_979 ();
 sg13g2_decap_8 FILLER_38_986 ();
 sg13g2_decap_8 FILLER_38_993 ();
 sg13g2_decap_8 FILLER_38_1000 ();
 sg13g2_decap_8 FILLER_38_1007 ();
 sg13g2_decap_8 FILLER_38_1014 ();
 sg13g2_decap_8 FILLER_38_1021 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_23 ();
 sg13g2_decap_4 FILLER_39_30 ();
 sg13g2_fill_2 FILLER_39_34 ();
 sg13g2_fill_2 FILLER_39_40 ();
 sg13g2_decap_4 FILLER_39_46 ();
 sg13g2_fill_1 FILLER_39_50 ();
 sg13g2_fill_1 FILLER_39_65 ();
 sg13g2_decap_8 FILLER_39_72 ();
 sg13g2_decap_8 FILLER_39_79 ();
 sg13g2_fill_2 FILLER_39_86 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_110 ();
 sg13g2_decap_4 FILLER_39_117 ();
 sg13g2_decap_8 FILLER_39_131 ();
 sg13g2_fill_2 FILLER_39_138 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_fill_1 FILLER_39_165 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_decap_4 FILLER_39_181 ();
 sg13g2_fill_1 FILLER_39_185 ();
 sg13g2_fill_2 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_238 ();
 sg13g2_decap_4 FILLER_39_245 ();
 sg13g2_fill_1 FILLER_39_249 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_2 FILLER_39_267 ();
 sg13g2_fill_1 FILLER_39_269 ();
 sg13g2_decap_8 FILLER_39_274 ();
 sg13g2_decap_4 FILLER_39_285 ();
 sg13g2_decap_4 FILLER_39_299 ();
 sg13g2_fill_2 FILLER_39_340 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_decap_4 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_414 ();
 sg13g2_fill_1 FILLER_39_416 ();
 sg13g2_fill_2 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_fill_1 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_446 ();
 sg13g2_decap_4 FILLER_39_453 ();
 sg13g2_fill_1 FILLER_39_457 ();
 sg13g2_decap_4 FILLER_39_468 ();
 sg13g2_fill_2 FILLER_39_472 ();
 sg13g2_decap_4 FILLER_39_496 ();
 sg13g2_decap_8 FILLER_39_527 ();
 sg13g2_decap_8 FILLER_39_534 ();
 sg13g2_decap_4 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_549 ();
 sg13g2_decap_8 FILLER_39_575 ();
 sg13g2_fill_1 FILLER_39_582 ();
 sg13g2_fill_2 FILLER_39_600 ();
 sg13g2_fill_1 FILLER_39_602 ();
 sg13g2_decap_4 FILLER_39_620 ();
 sg13g2_fill_1 FILLER_39_660 ();
 sg13g2_decap_8 FILLER_39_666 ();
 sg13g2_decap_8 FILLER_39_673 ();
 sg13g2_fill_1 FILLER_39_680 ();
 sg13g2_decap_4 FILLER_39_695 ();
 sg13g2_fill_1 FILLER_39_699 ();
 sg13g2_decap_8 FILLER_39_762 ();
 sg13g2_fill_2 FILLER_39_769 ();
 sg13g2_decap_4 FILLER_39_781 ();
 sg13g2_fill_2 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_fill_2 FILLER_39_868 ();
 sg13g2_fill_1 FILLER_39_870 ();
 sg13g2_decap_4 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_879 ();
 sg13g2_fill_1 FILLER_39_912 ();
 sg13g2_decap_8 FILLER_39_919 ();
 sg13g2_decap_8 FILLER_39_926 ();
 sg13g2_decap_4 FILLER_39_933 ();
 sg13g2_fill_1 FILLER_39_937 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1000 ();
 sg13g2_decap_8 FILLER_39_1007 ();
 sg13g2_decap_8 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1021 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_4 ();
 sg13g2_decap_4 FILLER_40_9 ();
 sg13g2_fill_2 FILLER_40_13 ();
 sg13g2_decap_8 FILLER_40_19 ();
 sg13g2_decap_4 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_decap_8 FILLER_40_76 ();
 sg13g2_decap_4 FILLER_40_83 ();
 sg13g2_fill_2 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_110 ();
 sg13g2_decap_8 FILLER_40_142 ();
 sg13g2_decap_4 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_153 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_fill_2 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_215 ();
 sg13g2_decap_8 FILLER_40_220 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_decap_4 FILLER_40_259 ();
 sg13g2_fill_2 FILLER_40_263 ();
 sg13g2_decap_4 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_fill_1 FILLER_40_336 ();
 sg13g2_fill_1 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_decap_4 FILLER_40_366 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_decap_4 FILLER_40_415 ();
 sg13g2_fill_1 FILLER_40_459 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_489 ();
 sg13g2_decap_4 FILLER_40_500 ();
 sg13g2_fill_1 FILLER_40_504 ();
 sg13g2_decap_4 FILLER_40_509 ();
 sg13g2_decap_8 FILLER_40_517 ();
 sg13g2_decap_8 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_531 ();
 sg13g2_fill_2 FILLER_40_538 ();
 sg13g2_decap_8 FILLER_40_566 ();
 sg13g2_fill_1 FILLER_40_573 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_594 ();
 sg13g2_fill_1 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_622 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_4 FILLER_40_658 ();
 sg13g2_decap_4 FILLER_40_698 ();
 sg13g2_decap_4 FILLER_40_732 ();
 sg13g2_decap_4 FILLER_40_775 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_fill_2 FILLER_40_828 ();
 sg13g2_fill_1 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_871 ();
 sg13g2_decap_4 FILLER_40_878 ();
 sg13g2_fill_2 FILLER_40_882 ();
 sg13g2_fill_1 FILLER_40_888 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_decap_4 FILLER_40_900 ();
 sg13g2_fill_2 FILLER_40_904 ();
 sg13g2_decap_4 FILLER_40_937 ();
 sg13g2_fill_1 FILLER_40_941 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_984 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_8 FILLER_40_998 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_fill_2 FILLER_40_1026 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_decap_8 FILLER_41_37 ();
 sg13g2_decap_8 FILLER_41_44 ();
 sg13g2_decap_4 FILLER_41_51 ();
 sg13g2_fill_1 FILLER_41_55 ();
 sg13g2_decap_4 FILLER_41_83 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_decap_8 FILLER_41_134 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_decap_8 FILLER_41_148 ();
 sg13g2_decap_4 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_decap_4 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_229 ();
 sg13g2_decap_4 FILLER_41_236 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_decap_4 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_260 ();
 sg13g2_decap_8 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_274 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_302 ();
 sg13g2_decap_8 FILLER_41_309 ();
 sg13g2_decap_4 FILLER_41_316 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_fill_2 FILLER_41_393 ();
 sg13g2_fill_1 FILLER_41_395 ();
 sg13g2_decap_8 FILLER_41_412 ();
 sg13g2_decap_4 FILLER_41_419 ();
 sg13g2_fill_2 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_41_435 ();
 sg13g2_decap_8 FILLER_41_442 ();
 sg13g2_decap_8 FILLER_41_449 ();
 sg13g2_decap_8 FILLER_41_456 ();
 sg13g2_fill_2 FILLER_41_463 ();
 sg13g2_decap_4 FILLER_41_469 ();
 sg13g2_fill_2 FILLER_41_473 ();
 sg13g2_decap_8 FILLER_41_479 ();
 sg13g2_decap_4 FILLER_41_486 ();
 sg13g2_decap_8 FILLER_41_530 ();
 sg13g2_fill_2 FILLER_41_537 ();
 sg13g2_decap_4 FILLER_41_567 ();
 sg13g2_fill_1 FILLER_41_583 ();
 sg13g2_decap_8 FILLER_41_601 ();
 sg13g2_decap_4 FILLER_41_608 ();
 sg13g2_fill_1 FILLER_41_617 ();
 sg13g2_decap_4 FILLER_41_623 ();
 sg13g2_fill_1 FILLER_41_627 ();
 sg13g2_decap_8 FILLER_41_632 ();
 sg13g2_decap_4 FILLER_41_639 ();
 sg13g2_fill_1 FILLER_41_643 ();
 sg13g2_decap_4 FILLER_41_662 ();
 sg13g2_fill_2 FILLER_41_666 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_fill_1 FILLER_41_679 ();
 sg13g2_decap_4 FILLER_41_684 ();
 sg13g2_decap_4 FILLER_41_728 ();
 sg13g2_fill_1 FILLER_41_732 ();
 sg13g2_decap_4 FILLER_41_760 ();
 sg13g2_fill_2 FILLER_41_794 ();
 sg13g2_fill_2 FILLER_41_855 ();
 sg13g2_fill_2 FILLER_41_884 ();
 sg13g2_fill_1 FILLER_41_886 ();
 sg13g2_decap_8 FILLER_41_919 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_decap_8 FILLER_41_933 ();
 sg13g2_fill_2 FILLER_41_940 ();
 sg13g2_fill_1 FILLER_41_942 ();
 sg13g2_decap_8 FILLER_41_951 ();
 sg13g2_decap_8 FILLER_41_958 ();
 sg13g2_decap_8 FILLER_41_965 ();
 sg13g2_decap_8 FILLER_41_972 ();
 sg13g2_decap_8 FILLER_41_979 ();
 sg13g2_decap_8 FILLER_41_986 ();
 sg13g2_decap_8 FILLER_41_993 ();
 sg13g2_decap_8 FILLER_41_1000 ();
 sg13g2_decap_8 FILLER_41_1007 ();
 sg13g2_decap_8 FILLER_41_1014 ();
 sg13g2_decap_8 FILLER_41_1021 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_11 ();
 sg13g2_fill_2 FILLER_42_17 ();
 sg13g2_fill_1 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_34 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_fill_2 FILLER_42_66 ();
 sg13g2_decap_8 FILLER_42_72 ();
 sg13g2_fill_2 FILLER_42_79 ();
 sg13g2_decap_8 FILLER_42_86 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_decap_4 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_156 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_187 ();
 sg13g2_decap_4 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_226 ();
 sg13g2_decap_4 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_324 ();
 sg13g2_decap_4 FILLER_42_331 ();
 sg13g2_decap_4 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_359 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_fill_2 FILLER_42_435 ();
 sg13g2_fill_1 FILLER_42_437 ();
 sg13g2_decap_4 FILLER_42_452 ();
 sg13g2_fill_2 FILLER_42_456 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_474 ();
 sg13g2_decap_4 FILLER_42_481 ();
 sg13g2_fill_1 FILLER_42_485 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_4 FILLER_42_504 ();
 sg13g2_fill_2 FILLER_42_512 ();
 sg13g2_fill_1 FILLER_42_514 ();
 sg13g2_decap_8 FILLER_42_519 ();
 sg13g2_decap_8 FILLER_42_526 ();
 sg13g2_decap_4 FILLER_42_533 ();
 sg13g2_fill_1 FILLER_42_537 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_fill_2 FILLER_42_573 ();
 sg13g2_decap_8 FILLER_42_593 ();
 sg13g2_decap_4 FILLER_42_600 ();
 sg13g2_fill_1 FILLER_42_604 ();
 sg13g2_decap_4 FILLER_42_627 ();
 sg13g2_fill_1 FILLER_42_631 ();
 sg13g2_fill_1 FILLER_42_649 ();
 sg13g2_decap_4 FILLER_42_654 ();
 sg13g2_fill_2 FILLER_42_743 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_4 FILLER_42_789 ();
 sg13g2_fill_2 FILLER_42_793 ();
 sg13g2_fill_1 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_891 ();
 sg13g2_decap_8 FILLER_42_902 ();
 sg13g2_decap_8 FILLER_42_909 ();
 sg13g2_decap_8 FILLER_42_916 ();
 sg13g2_decap_8 FILLER_42_923 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_8 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_8 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_54 ();
 sg13g2_decap_8 FILLER_43_61 ();
 sg13g2_fill_2 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_fill_2 FILLER_43_184 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_fill_1 FILLER_43_240 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_decap_4 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_299 ();
 sg13g2_fill_2 FILLER_43_306 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_decap_4 FILLER_43_399 ();
 sg13g2_decap_4 FILLER_43_430 ();
 sg13g2_decap_8 FILLER_43_461 ();
 sg13g2_decap_8 FILLER_43_468 ();
 sg13g2_fill_1 FILLER_43_493 ();
 sg13g2_decap_8 FILLER_43_498 ();
 sg13g2_fill_2 FILLER_43_505 ();
 sg13g2_decap_8 FILLER_43_534 ();
 sg13g2_decap_4 FILLER_43_541 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_fill_2 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_decap_8 FILLER_43_597 ();
 sg13g2_fill_1 FILLER_43_604 ();
 sg13g2_fill_1 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_619 ();
 sg13g2_decap_4 FILLER_43_626 ();
 sg13g2_fill_2 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_decap_8 FILLER_43_666 ();
 sg13g2_decap_8 FILLER_43_673 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_4 FILLER_43_691 ();
 sg13g2_decap_4 FILLER_43_699 ();
 sg13g2_fill_1 FILLER_43_703 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_fill_2 FILLER_43_781 ();
 sg13g2_fill_1 FILLER_43_783 ();
 sg13g2_fill_1 FILLER_43_794 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_fill_2 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_4 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_893 ();
 sg13g2_decap_8 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_907 ();
 sg13g2_decap_8 FILLER_43_914 ();
 sg13g2_decap_8 FILLER_43_921 ();
 sg13g2_decap_8 FILLER_43_928 ();
 sg13g2_decap_8 FILLER_43_935 ();
 sg13g2_decap_8 FILLER_43_942 ();
 sg13g2_decap_8 FILLER_43_949 ();
 sg13g2_decap_8 FILLER_43_956 ();
 sg13g2_decap_8 FILLER_43_963 ();
 sg13g2_decap_8 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_977 ();
 sg13g2_decap_8 FILLER_43_984 ();
 sg13g2_decap_8 FILLER_43_991 ();
 sg13g2_decap_8 FILLER_43_998 ();
 sg13g2_decap_8 FILLER_43_1005 ();
 sg13g2_decap_8 FILLER_43_1012 ();
 sg13g2_decap_8 FILLER_43_1019 ();
 sg13g2_fill_2 FILLER_43_1026 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_42 ();
 sg13g2_decap_4 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_decap_4 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_159 ();
 sg13g2_decap_8 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_fill_2 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_196 ();
 sg13g2_decap_4 FILLER_44_202 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_fill_2 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_214 ();
 sg13g2_fill_1 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_fill_2 FILLER_44_259 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_4 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_fill_2 FILLER_44_294 ();
 sg13g2_decap_4 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_310 ();
 sg13g2_fill_2 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_317 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_decap_8 FILLER_44_365 ();
 sg13g2_decap_4 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_376 ();
 sg13g2_decap_4 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_fill_1 FILLER_44_407 ();
 sg13g2_fill_2 FILLER_44_412 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_4 FILLER_44_431 ();
 sg13g2_fill_1 FILLER_44_435 ();
 sg13g2_decap_8 FILLER_44_450 ();
 sg13g2_decap_4 FILLER_44_457 ();
 sg13g2_decap_8 FILLER_44_502 ();
 sg13g2_fill_2 FILLER_44_509 ();
 sg13g2_fill_1 FILLER_44_511 ();
 sg13g2_fill_1 FILLER_44_516 ();
 sg13g2_decap_8 FILLER_44_521 ();
 sg13g2_decap_8 FILLER_44_528 ();
 sg13g2_decap_8 FILLER_44_535 ();
 sg13g2_decap_4 FILLER_44_542 ();
 sg13g2_fill_2 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_552 ();
 sg13g2_decap_8 FILLER_44_559 ();
 sg13g2_decap_8 FILLER_44_566 ();
 sg13g2_decap_4 FILLER_44_573 ();
 sg13g2_fill_1 FILLER_44_577 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_4 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_4 FILLER_44_641 ();
 sg13g2_fill_2 FILLER_44_645 ();
 sg13g2_fill_2 FILLER_44_678 ();
 sg13g2_fill_1 FILLER_44_680 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_fill_2 FILLER_44_746 ();
 sg13g2_fill_1 FILLER_44_748 ();
 sg13g2_decap_4 FILLER_44_759 ();
 sg13g2_fill_2 FILLER_44_763 ();
 sg13g2_fill_1 FILLER_44_792 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_4 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_883 ();
 sg13g2_decap_8 FILLER_44_890 ();
 sg13g2_decap_8 FILLER_44_897 ();
 sg13g2_decap_8 FILLER_44_904 ();
 sg13g2_decap_8 FILLER_44_911 ();
 sg13g2_decap_8 FILLER_44_918 ();
 sg13g2_decap_8 FILLER_44_925 ();
 sg13g2_decap_8 FILLER_44_932 ();
 sg13g2_decap_8 FILLER_44_939 ();
 sg13g2_decap_8 FILLER_44_946 ();
 sg13g2_decap_8 FILLER_44_953 ();
 sg13g2_decap_8 FILLER_44_960 ();
 sg13g2_decap_8 FILLER_44_967 ();
 sg13g2_decap_8 FILLER_44_974 ();
 sg13g2_decap_8 FILLER_44_981 ();
 sg13g2_decap_8 FILLER_44_988 ();
 sg13g2_decap_8 FILLER_44_995 ();
 sg13g2_decap_8 FILLER_44_1002 ();
 sg13g2_decap_8 FILLER_44_1009 ();
 sg13g2_decap_8 FILLER_44_1016 ();
 sg13g2_decap_4 FILLER_44_1023 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_decap_4 FILLER_45_22 ();
 sg13g2_fill_2 FILLER_45_26 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_fill_1 FILLER_45_34 ();
 sg13g2_decap_8 FILLER_45_45 ();
 sg13g2_decap_8 FILLER_45_52 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_73 ();
 sg13g2_decap_8 FILLER_45_80 ();
 sg13g2_decap_8 FILLER_45_87 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_fill_2 FILLER_45_170 ();
 sg13g2_decap_4 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_fill_2 FILLER_45_337 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_fill_1 FILLER_45_397 ();
 sg13g2_fill_1 FILLER_45_435 ();
 sg13g2_decap_8 FILLER_45_467 ();
 sg13g2_decap_4 FILLER_45_474 ();
 sg13g2_fill_2 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_484 ();
 sg13g2_decap_4 FILLER_45_491 ();
 sg13g2_fill_2 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_507 ();
 sg13g2_decap_8 FILLER_45_535 ();
 sg13g2_fill_1 FILLER_45_542 ();
 sg13g2_fill_2 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_573 ();
 sg13g2_decap_8 FILLER_45_618 ();
 sg13g2_decap_8 FILLER_45_625 ();
 sg13g2_decap_4 FILLER_45_632 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_752 ();
 sg13g2_fill_1 FILLER_45_759 ();
 sg13g2_decap_4 FILLER_45_804 ();
 sg13g2_decap_4 FILLER_45_867 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_decap_8 FILLER_45_887 ();
 sg13g2_decap_8 FILLER_45_894 ();
 sg13g2_decap_8 FILLER_45_901 ();
 sg13g2_decap_8 FILLER_45_908 ();
 sg13g2_decap_8 FILLER_45_915 ();
 sg13g2_decap_8 FILLER_45_922 ();
 sg13g2_decap_8 FILLER_45_929 ();
 sg13g2_decap_8 FILLER_45_936 ();
 sg13g2_decap_8 FILLER_45_943 ();
 sg13g2_decap_8 FILLER_45_950 ();
 sg13g2_decap_8 FILLER_45_957 ();
 sg13g2_decap_8 FILLER_45_964 ();
 sg13g2_decap_8 FILLER_45_971 ();
 sg13g2_decap_8 FILLER_45_978 ();
 sg13g2_decap_8 FILLER_45_985 ();
 sg13g2_decap_8 FILLER_45_992 ();
 sg13g2_decap_8 FILLER_45_999 ();
 sg13g2_decap_8 FILLER_45_1006 ();
 sg13g2_decap_8 FILLER_45_1013 ();
 sg13g2_decap_4 FILLER_45_1020 ();
 sg13g2_fill_1 FILLER_45_1024 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_decap_4 FILLER_46_60 ();
 sg13g2_fill_2 FILLER_46_64 ();
 sg13g2_fill_2 FILLER_46_74 ();
 sg13g2_fill_1 FILLER_46_76 ();
 sg13g2_decap_4 FILLER_46_95 ();
 sg13g2_fill_1 FILLER_46_99 ();
 sg13g2_fill_2 FILLER_46_121 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_decap_4 FILLER_46_181 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_decap_4 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_decap_4 FILLER_46_251 ();
 sg13g2_decap_8 FILLER_46_267 ();
 sg13g2_decap_4 FILLER_46_274 ();
 sg13g2_fill_1 FILLER_46_278 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_4 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_309 ();
 sg13g2_fill_2 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_decap_4 FILLER_46_323 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_fill_2 FILLER_46_339 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_decap_8 FILLER_46_369 ();
 sg13g2_fill_2 FILLER_46_376 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_46_425 ();
 sg13g2_decap_8 FILLER_46_432 ();
 sg13g2_decap_4 FILLER_46_439 ();
 sg13g2_fill_1 FILLER_46_443 ();
 sg13g2_decap_4 FILLER_46_456 ();
 sg13g2_fill_2 FILLER_46_464 ();
 sg13g2_fill_1 FILLER_46_466 ();
 sg13g2_decap_8 FILLER_46_477 ();
 sg13g2_fill_2 FILLER_46_493 ();
 sg13g2_fill_1 FILLER_46_495 ();
 sg13g2_decap_8 FILLER_46_500 ();
 sg13g2_decap_4 FILLER_46_507 ();
 sg13g2_fill_2 FILLER_46_511 ();
 sg13g2_fill_1 FILLER_46_517 ();
 sg13g2_decap_8 FILLER_46_522 ();
 sg13g2_decap_8 FILLER_46_529 ();
 sg13g2_decap_8 FILLER_46_536 ();
 sg13g2_decap_4 FILLER_46_543 ();
 sg13g2_fill_1 FILLER_46_547 ();
 sg13g2_fill_1 FILLER_46_576 ();
 sg13g2_decap_4 FILLER_46_590 ();
 sg13g2_fill_1 FILLER_46_594 ();
 sg13g2_fill_1 FILLER_46_622 ();
 sg13g2_decap_4 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_659 ();
 sg13g2_decap_4 FILLER_46_694 ();
 sg13g2_fill_2 FILLER_46_698 ();
 sg13g2_fill_1 FILLER_46_736 ();
 sg13g2_fill_2 FILLER_46_749 ();
 sg13g2_fill_1 FILLER_46_751 ();
 sg13g2_decap_4 FILLER_46_761 ();
 sg13g2_fill_1 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_decap_8 FILLER_46_782 ();
 sg13g2_decap_8 FILLER_46_789 ();
 sg13g2_decap_8 FILLER_46_796 ();
 sg13g2_decap_8 FILLER_46_803 ();
 sg13g2_decap_8 FILLER_46_810 ();
 sg13g2_decap_4 FILLER_46_817 ();
 sg13g2_fill_2 FILLER_46_821 ();
 sg13g2_fill_1 FILLER_46_832 ();
 sg13g2_decap_4 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_846 ();
 sg13g2_decap_4 FILLER_46_851 ();
 sg13g2_fill_1 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_46_865 ();
 sg13g2_decap_8 FILLER_46_872 ();
 sg13g2_decap_8 FILLER_46_879 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_decap_8 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_900 ();
 sg13g2_decap_8 FILLER_46_907 ();
 sg13g2_decap_8 FILLER_46_914 ();
 sg13g2_decap_8 FILLER_46_921 ();
 sg13g2_decap_8 FILLER_46_928 ();
 sg13g2_decap_8 FILLER_46_935 ();
 sg13g2_decap_8 FILLER_46_942 ();
 sg13g2_decap_8 FILLER_46_949 ();
 sg13g2_decap_8 FILLER_46_956 ();
 sg13g2_decap_8 FILLER_46_963 ();
 sg13g2_decap_8 FILLER_46_970 ();
 sg13g2_decap_8 FILLER_46_977 ();
 sg13g2_decap_8 FILLER_46_984 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_998 ();
 sg13g2_decap_8 FILLER_46_1005 ();
 sg13g2_decap_8 FILLER_46_1012 ();
 sg13g2_decap_8 FILLER_46_1019 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_fill_2 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_147 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_162 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_4 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_189 ();
 sg13g2_decap_4 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_229 ();
 sg13g2_fill_1 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_decap_8 FILLER_47_334 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_4 FILLER_47_379 ();
 sg13g2_fill_2 FILLER_47_387 ();
 sg13g2_fill_1 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_decap_8 FILLER_47_425 ();
 sg13g2_decap_4 FILLER_47_432 ();
 sg13g2_fill_2 FILLER_47_446 ();
 sg13g2_fill_1 FILLER_47_448 ();
 sg13g2_decap_4 FILLER_47_489 ();
 sg13g2_fill_1 FILLER_47_493 ();
 sg13g2_fill_1 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_557 ();
 sg13g2_decap_8 FILLER_47_564 ();
 sg13g2_decap_8 FILLER_47_571 ();
 sg13g2_decap_8 FILLER_47_578 ();
 sg13g2_decap_8 FILLER_47_585 ();
 sg13g2_decap_8 FILLER_47_592 ();
 sg13g2_fill_1 FILLER_47_599 ();
 sg13g2_decap_8 FILLER_47_604 ();
 sg13g2_decap_8 FILLER_47_611 ();
 sg13g2_decap_8 FILLER_47_618 ();
 sg13g2_fill_2 FILLER_47_652 ();
 sg13g2_decap_8 FILLER_47_663 ();
 sg13g2_fill_2 FILLER_47_670 ();
 sg13g2_fill_2 FILLER_47_709 ();
 sg13g2_fill_1 FILLER_47_711 ();
 sg13g2_fill_1 FILLER_47_725 ();
 sg13g2_fill_2 FILLER_47_795 ();
 sg13g2_fill_1 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_decap_8 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_871 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_8 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_983 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_61 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_decap_4 FILLER_48_75 ();
 sg13g2_decap_8 FILLER_48_87 ();
 sg13g2_decap_8 FILLER_48_94 ();
 sg13g2_decap_8 FILLER_48_101 ();
 sg13g2_decap_8 FILLER_48_108 ();
 sg13g2_fill_2 FILLER_48_115 ();
 sg13g2_decap_8 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_decap_4 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_210 ();
 sg13g2_decap_4 FILLER_48_239 ();
 sg13g2_decap_4 FILLER_48_307 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_decap_8 FILLER_48_358 ();
 sg13g2_decap_8 FILLER_48_365 ();
 sg13g2_decap_8 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_decap_8 FILLER_48_386 ();
 sg13g2_decap_8 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_409 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_466 ();
 sg13g2_decap_4 FILLER_48_471 ();
 sg13g2_decap_8 FILLER_48_479 ();
 sg13g2_decap_8 FILLER_48_486 ();
 sg13g2_decap_8 FILLER_48_493 ();
 sg13g2_decap_8 FILLER_48_500 ();
 sg13g2_fill_2 FILLER_48_507 ();
 sg13g2_fill_1 FILLER_48_509 ();
 sg13g2_fill_2 FILLER_48_514 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_527 ();
 sg13g2_decap_8 FILLER_48_534 ();
 sg13g2_decap_8 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_548 ();
 sg13g2_decap_8 FILLER_48_555 ();
 sg13g2_decap_8 FILLER_48_562 ();
 sg13g2_decap_8 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_decap_8 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_597 ();
 sg13g2_decap_8 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_decap_4 FILLER_48_625 ();
 sg13g2_fill_1 FILLER_48_629 ();
 sg13g2_decap_8 FILLER_48_634 ();
 sg13g2_decap_8 FILLER_48_641 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_decap_8 FILLER_48_655 ();
 sg13g2_fill_2 FILLER_48_690 ();
 sg13g2_fill_2 FILLER_48_705 ();
 sg13g2_fill_1 FILLER_48_707 ();
 sg13g2_fill_1 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_fill_2 FILLER_48_754 ();
 sg13g2_decap_4 FILLER_48_792 ();
 sg13g2_fill_2 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_867 ();
 sg13g2_decap_8 FILLER_48_874 ();
 sg13g2_decap_8 FILLER_48_881 ();
 sg13g2_decap_8 FILLER_48_888 ();
 sg13g2_decap_8 FILLER_48_895 ();
 sg13g2_decap_8 FILLER_48_902 ();
 sg13g2_decap_8 FILLER_48_909 ();
 sg13g2_decap_8 FILLER_48_916 ();
 sg13g2_decap_8 FILLER_48_923 ();
 sg13g2_decap_8 FILLER_48_930 ();
 sg13g2_decap_8 FILLER_48_937 ();
 sg13g2_decap_8 FILLER_48_944 ();
 sg13g2_decap_8 FILLER_48_951 ();
 sg13g2_decap_8 FILLER_48_958 ();
 sg13g2_decap_8 FILLER_48_965 ();
 sg13g2_decap_8 FILLER_48_972 ();
 sg13g2_decap_8 FILLER_48_979 ();
 sg13g2_decap_8 FILLER_48_986 ();
 sg13g2_decap_8 FILLER_48_993 ();
 sg13g2_decap_8 FILLER_48_1000 ();
 sg13g2_decap_8 FILLER_48_1007 ();
 sg13g2_decap_8 FILLER_48_1014 ();
 sg13g2_decap_8 FILLER_48_1021 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_4 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_127 ();
 sg13g2_decap_8 FILLER_49_134 ();
 sg13g2_decap_8 FILLER_49_141 ();
 sg13g2_decap_8 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_decap_8 FILLER_49_160 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_8 FILLER_49_174 ();
 sg13g2_fill_2 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_decap_8 FILLER_49_188 ();
 sg13g2_decap_8 FILLER_49_195 ();
 sg13g2_decap_8 FILLER_49_202 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_decap_4 FILLER_49_224 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_247 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_fill_2 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_272 ();
 sg13g2_decap_4 FILLER_49_279 ();
 sg13g2_fill_2 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_decap_8 FILLER_49_296 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_338 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_8 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_387 ();
 sg13g2_decap_8 FILLER_49_394 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_decap_8 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_426 ();
 sg13g2_decap_8 FILLER_49_433 ();
 sg13g2_decap_4 FILLER_49_440 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_fill_1 FILLER_49_651 ();
 sg13g2_fill_2 FILLER_49_723 ();
 sg13g2_decap_8 FILLER_49_730 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_8 FILLER_49_744 ();
 sg13g2_decap_8 FILLER_49_751 ();
 sg13g2_fill_2 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_fill_2 FILLER_49_779 ();
 sg13g2_fill_1 FILLER_49_781 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_834 ();
 sg13g2_decap_8 FILLER_49_841 ();
 sg13g2_decap_8 FILLER_49_848 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_decap_8 FILLER_49_862 ();
 sg13g2_decap_8 FILLER_49_869 ();
 sg13g2_decap_8 FILLER_49_876 ();
 sg13g2_decap_8 FILLER_49_883 ();
 sg13g2_decap_8 FILLER_49_890 ();
 sg13g2_decap_8 FILLER_49_897 ();
 sg13g2_decap_8 FILLER_49_904 ();
 sg13g2_decap_8 FILLER_49_911 ();
 sg13g2_decap_8 FILLER_49_918 ();
 sg13g2_decap_8 FILLER_49_925 ();
 sg13g2_decap_8 FILLER_49_932 ();
 sg13g2_decap_8 FILLER_49_939 ();
 sg13g2_decap_8 FILLER_49_946 ();
 sg13g2_decap_8 FILLER_49_953 ();
 sg13g2_decap_8 FILLER_49_960 ();
 sg13g2_decap_8 FILLER_49_967 ();
 sg13g2_decap_8 FILLER_49_974 ();
 sg13g2_decap_8 FILLER_49_981 ();
 sg13g2_decap_8 FILLER_49_988 ();
 sg13g2_decap_8 FILLER_49_995 ();
 sg13g2_decap_8 FILLER_49_1002 ();
 sg13g2_decap_8 FILLER_49_1009 ();
 sg13g2_decap_8 FILLER_49_1016 ();
 sg13g2_decap_4 FILLER_49_1023 ();
 sg13g2_fill_2 FILLER_49_1027 ();
 assign uio_oe[0] = net21;
 assign uio_oe[1] = net22;
 assign uio_oe[2] = net23;
 assign uio_oe[3] = net24;
 assign uio_oe[4] = net25;
 assign uio_oe[5] = net26;
 assign uio_oe[6] = net27;
 assign uio_oe[7] = net28;
 assign uio_out[1] = net29;
 assign uio_out[5] = net30;
endmodule
