* NGSPICE file created from heichips25_bagel.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

.subckt heichips25_bagel VGND VPWR clk ena rst_n tmds_b tmds_clk tmds_g tmds_r ui_in[0]
+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1]
+ uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_28_907 VPWR VGND sg13g2_decap_8
X_3155_ _0919_ _0925_ _0926_ _0321_ VPWR VGND sg13g2_nor3_1
XFILLER_39_299 VPWR VGND sg13g2_decap_4
X_3086_ _0865_ _0875_ _0876_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_439 VPWR VGND sg13g2_fill_1
XFILLER_36_940 VPWR VGND sg13g2_fill_1
X_4864__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_35_483 VPWR VGND sg13g2_decap_4
X_3988_ _1712_ _1713_ _1714_ VPWR VGND sg13g2_nor2_1
X_2939_ _0797_ videogen.fancy_shader.video_x\[3\] _0795_ VPWR VGND sg13g2_nand2_1
XFILLER_22_199 VPWR VGND sg13g2_decap_8
X_4609_ net690 net744 _0162_ VPWR VGND sg13g2_nor2_1
XFILLER_2_538 VPWR VGND sg13g2_fill_1
XFILLER_18_439 VPWR VGND sg13g2_decap_8
X_4982__269 VPWR VGND net269 sg13g2_tiehi
XFILLER_26_30 VPWR VGND sg13g2_decap_4
XFILLER_27_940 VPWR VGND sg13g2_decap_8
XFILLER_26_472 VPWR VGND sg13g2_fill_1
XFILLER_42_965 VPWR VGND sg13g2_decap_8
XFILLER_41_442 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk_regs clknet_0_clk_regs clknet_3_6__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_41_486 VPWR VGND sg13g2_decap_4
XFILLER_13_199 VPWR VGND sg13g2_fill_1
XFILLER_3_56 VPWR VGND sg13g2_decap_4
XFILLER_3_34 VPWR VGND sg13g2_fill_2
XFILLER_1_560 VPWR VGND sg13g2_fill_1
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_37_748 VPWR VGND sg13g2_decap_8
XFILLER_37_737 VPWR VGND sg13g2_fill_1
XFILLER_37_726 VPWR VGND sg13g2_decap_8
XFILLER_18_973 VPWR VGND sg13g2_decap_8
X_4960_ net379 VGND VPWR _0507_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\]
+ _0155_ sg13g2_dfrbpq_1
XFILLER_33_910 VPWR VGND sg13g2_fill_1
X_3911_ _1637_ _1124_ _1636_ VPWR VGND sg13g2_xnor2_1
X_4891_ net214 VGND VPWR _0442_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\]
+ _0099_ sg13g2_dfrbpq_1
XFILLER_33_965 VPWR VGND sg13g2_decap_8
X_3842_ net622 VPWR _1571_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\]
+ net580 sg13g2_o21ai_1
X_4785__32 VPWR VGND net32 sg13g2_tiehi
X_3773_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\] net553 _1503_ VPWR
+ VGND sg13g2_nor2_1
X_2724_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\] net780 _0744_ _0519_
+ VPWR VGND sg13g2_mux2_1
X_2655_ _0730_ _0698_ _0713_ VPWR VGND sg13g2_nand2_2
X_2586_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\] net752 _0700_ _0631_
+ VPWR VGND sg13g2_mux2_1
X_4325_ net601 tmds_green.n126 _2021_ VPWR VGND sg13g2_nor2_1
X_4256_ VGND VPWR _1940_ _1959_ _1962_ _1961_ sg13g2_a21oi_1
X_3207_ net751 _0959_ _0960_ _0347_ VPWR VGND sg13g2_nor3_1
X_4187_ _1619_ _1720_ _1351_ _1907_ VPWR VGND sg13g2_nand3_1
X_3138_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\]
+ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0913_ VPWR VGND sg13g2_nor3_1
XFILLER_28_748 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
X_3069_ tmds_red.n132 tmds_red.n114 _0859_ VPWR VGND sg13g2_xor2_1
XFILLER_24_932 VPWR VGND sg13g2_decap_8
XFILLER_23_442 VPWR VGND sg13g2_decap_8
XFILLER_3_869 VPWR VGND sg13g2_decap_8
Xfanout650 clk_video net650 VPWR VGND sg13g2_buf_8
Xfanout672 net673 net672 VPWR VGND sg13g2_buf_2
Xfanout694 clockdiv.q2temp net694 VPWR VGND sg13g2_buf_8
Xfanout683 net694 net683 VPWR VGND sg13g2_buf_8
Xfanout661 net663 net661 VPWR VGND sg13g2_buf_8
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_19_726 VPWR VGND sg13g2_decap_4
XFILLER_37_73 VPWR VGND sg13g2_decap_8
XFILLER_18_258 VPWR VGND sg13g2_decap_4
XFILLER_42_762 VPWR VGND sg13g2_decap_8
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_30_902 VPWR VGND sg13g2_decap_8
XFILLER_30_979 VPWR VGND sg13g2_decap_8
X_5090_ net801 VGND VPWR serialize.n428\[5\] serialize.n414\[3\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4110_ _1806_ _1826_ _1829_ _1833_ VPWR VGND sg13g2_nor3_1
X_4041_ VGND VPWR _1764_ _1757_ _1749_ sg13g2_or2_1
XFILLER_37_512 VPWR VGND sg13g2_fill_2
XFILLER_49_394 VPWR VGND sg13g2_decap_8
XFILLER_37_545 VPWR VGND sg13g2_decap_4
X_4943_ net57 VGND VPWR _0490_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\]
+ _0147_ sg13g2_dfrbpq_1
XFILLER_21_902 VPWR VGND sg13g2_fill_1
X_4874_ net247 VGND VPWR _0425_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\]
+ _0082_ sg13g2_dfrbpq_1
XFILLER_21_957 VPWR VGND sg13g2_decap_8
XFILLER_32_272 VPWR VGND sg13g2_decap_4
XFILLER_32_283 VPWR VGND sg13g2_decap_4
X_3825_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\] net555 _1554_ VPWR
+ VGND sg13g2_nor2_1
X_3756_ net615 VPWR _1486_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\]
+ net561 sg13g2_o21ai_1
X_2707_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\] _0741_ _0533_
+ VPWR VGND sg13g2_mux2_1
X_3687_ net596 VPWR _1417_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\]
+ net560 sg13g2_o21ai_1
X_2638_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\] net755 _0724_ _0585_
+ VPWR VGND sg13g2_mux2_1
X_4716__151 VPWR VGND net151 sg13g2_tiehi
XFILLER_0_828 VPWR VGND sg13g2_decap_8
X_2569_ _0684_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _0681_ VPWR VGND
+ sg13g2_xnor2_1
X_4308_ tmds_blue.n132 net605 _2008_ VPWR VGND sg13g2_xor2_1
X_4239_ VPWR _1946_ _1945_ VGND sg13g2_inv_1
XFILLER_24_740 VPWR VGND sg13g2_decap_8
XFILLER_12_946 VPWR VGND sg13g2_decap_8
XFILLER_23_20 VPWR VGND sg13g2_fill_1
XFILLER_24_784 VPWR VGND sg13g2_decap_8
XFILLER_11_445 VPWR VGND sg13g2_decap_8
XFILLER_3_677 VPWR VGND sg13g2_decap_8
XFILLER_2_132 VPWR VGND sg13g2_decap_8
X_4988__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_48_61 VPWR VGND sg13g2_decap_8
XFILLER_48_94 VPWR VGND sg13g2_decap_8
XFILLER_17_9 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_fill_1
XFILLER_0_79 VPWR VGND sg13g2_fill_1
XFILLER_30_710 VPWR VGND sg13g2_decap_8
XFILLER_9_66 VPWR VGND sg13g2_fill_1
X_3610_ _1336_ _1337_ _1338_ _1339_ _1340_ VPWR VGND sg13g2_nor4_1
XFILLER_30_787 VPWR VGND sg13g2_fill_2
X_4590_ net687 net738 _0143_ VPWR VGND sg13g2_nor2_1
X_3541_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\] net549 _1271_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_7_961 VPWR VGND sg13g2_decap_8
X_3472_ _1202_ _1066_ _1200_ VPWR VGND sg13g2_nand2_1
X_5073_ net122 VGND VPWR _0620_ tmds_green.dc_balancing_reg\[2\] net648 sg13g2_dfrbpq_1
X_4024_ _1739_ VPWR _1747_ VGND _1736_ _1742_ sg13g2_o21ai_1
X_4926_ net120 VGND VPWR _0477_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\]
+ _0134_ sg13g2_dfrbpq_1
X_4857_ net284 VGND VPWR _0408_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\]
+ _0065_ sg13g2_dfrbpq_1
X_3808_ _1534_ _1535_ _1536_ _1537_ _1538_ VPWR VGND sg13g2_nor4_1
X_4800__374 VPWR VGND net374 sg13g2_tiehi
X_4788_ net398 VGND VPWR _0339_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\]
+ _0039_ sg13g2_dfrbpq_1
X_3739_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\] net574 _1469_ VPWR
+ VGND sg13g2_nor2_1
Xheichips25_bagel_24 VPWR VGND uio_oe[3] sg13g2_tielo
XFILLER_0_625 VPWR VGND sg13g2_fill_2
XFILLER_48_618 VPWR VGND sg13g2_decap_8
XFILLER_48_629 VPWR VGND sg13g2_fill_1
XFILLER_29_810 VPWR VGND sg13g2_decap_4
XFILLER_28_353 VPWR VGND sg13g2_fill_1
XFILLER_43_312 VPWR VGND sg13g2_fill_1
XFILLER_11_220 VPWR VGND sg13g2_decap_4
XFILLER_12_754 VPWR VGND sg13g2_decap_8
XFILLER_24_592 VPWR VGND sg13g2_decap_8
XFILLER_11_275 VPWR VGND sg13g2_fill_1
XFILLER_8_758 VPWR VGND sg13g2_decap_4
XFILLER_4_964 VPWR VGND sg13g2_decap_8
X_5062__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_34_301 VPWR VGND sg13g2_fill_1
XFILLER_35_879 VPWR VGND sg13g2_decap_4
X_2972_ net600 VPWR _0820_ VGND _0813_ _0818_ sg13g2_o21ai_1
X_4711_ net253 VGND VPWR _0263_ tmds_green.dc_balancing_reg\[0\] net648 sg13g2_dfrbpq_1
XFILLER_30_540 VPWR VGND sg13g2_decap_4
X_4642_ net664 net715 _0195_ VPWR VGND sg13g2_nor2_1
X_4573_ net676 net728 _0126_ VPWR VGND sg13g2_nor2_1
X_3524_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\] net560 _1254_ VPWR
+ VGND sg13g2_nor2_1
X_3455_ _1147_ VPWR _1185_ VGND _1156_ _1183_ sg13g2_o21ai_1
X_3386_ VGND VPWR _1080_ _1082_ _1116_ _1081_ sg13g2_a21oi_1
X_4713__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_29_106 VPWR VGND sg13g2_decap_8
X_5125_ net798 VGND VPWR serialize.n427\[9\] serialize.n411\[7\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5056_ net361 VGND VPWR _0603_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\]
+ _0251_ sg13g2_dfrbpq_1
X_4007_ _1730_ _1076_ _1729_ VPWR VGND sg13g2_nand2_1
XFILLER_26_824 VPWR VGND sg13g2_fill_1
XFILLER_25_323 VPWR VGND sg13g2_fill_1
XFILLER_26_857 VPWR VGND sg13g2_fill_1
XFILLER_38_1007 VPWR VGND sg13g2_decap_8
XFILLER_26_868 VPWR VGND sg13g2_fill_2
XFILLER_40_359 VPWR VGND sg13g2_decap_8
X_4909_ net178 VGND VPWR _0460_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\]
+ _0117_ sg13g2_dfrbpq_1
X_4978__285 VPWR VGND net285 sg13g2_tiehi
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_4_216 VPWR VGND sg13g2_decap_8
XFILLER_20_43 VPWR VGND sg13g2_fill_1
XFILLER_20_76 VPWR VGND sg13g2_decap_4
XFILLER_1_923 VPWR VGND sg13g2_decap_8
Xhold41 _0004_ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold30 serialize.n411\[4\] VPWR VGND net435 sg13g2_dlygate4sd3_1
XFILLER_48_437 VPWR VGND sg13g2_fill_2
XFILLER_29_85 VPWR VGND sg13g2_decap_8
XFILLER_35_109 VPWR VGND sg13g2_fill_1
XFILLER_28_172 VPWR VGND sg13g2_fill_1
XFILLER_45_73 VPWR VGND sg13g2_decap_8
XFILLER_16_367 VPWR VGND sg13g2_fill_2
XFILLER_44_698 VPWR VGND sg13g2_decap_8
X_4992__227 VPWR VGND net227 sg13g2_tiehi
XFILLER_40_882 VPWR VGND sg13g2_fill_2
XFILLER_40_871 VPWR VGND sg13g2_decap_8
XFILLER_40_893 VPWR VGND sg13g2_decap_8
XFILLER_6_34 VPWR VGND sg13g2_fill_1
X_3240_ _0981_ _0982_ _0358_ VPWR VGND sg13g2_nor2_1
XFILLER_39_404 VPWR VGND sg13g2_decap_4
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
X_3171_ net621 _0935_ _0938_ VPWR VGND sg13g2_and2_1
XFILLER_48_993 VPWR VGND sg13g2_decap_8
XFILLER_23_805 VPWR VGND sg13g2_decap_8
XFILLER_16_890 VPWR VGND sg13g2_fill_1
X_2955_ _0792_ VPWR _0812_ VGND videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ _0807_ sg13g2_o21ai_1
X_2886_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\] net782 _0781_ _0342_
+ VPWR VGND sg13g2_mux2_1
X_4625_ net689 net741 _0178_ VPWR VGND sg13g2_nor2_1
X_4556_ net682 net733 _0109_ VPWR VGND sg13g2_nor2_1
X_3507_ VGND VPWR _1237_ _1231_ _1176_ sg13g2_or2_1
X_4487_ net685 net736 _0040_ VPWR VGND sg13g2_nor2_1
X_3438_ _1153_ VPWR _1168_ VGND _1152_ _1167_ sg13g2_o21ai_1
X_3369_ _1099_ _1097_ _1098_ VPWR VGND sg13g2_xnor2_1
X_5108_ net800 VGND VPWR serialize.n429\[5\] serialize.n417\[3\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_39_993 VPWR VGND sg13g2_decap_8
X_5039_ net229 VGND VPWR _0586_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\]
+ _0234_ sg13g2_dfrbpq_1
XFILLER_26_643 VPWR VGND sg13g2_decap_8
XFILLER_14_849 VPWR VGND sg13g2_decap_4
XFILLER_15_21 VPWR VGND sg13g2_fill_1
XFILLER_15_65 VPWR VGND sg13g2_fill_1
XFILLER_41_679 VPWR VGND sg13g2_fill_1
Xclkbuf_3_5__f_clk_regs clknet_0_clk_regs clknet_3_5__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_15_76 VPWR VGND sg13g2_fill_2
XFILLER_15_98 VPWR VGND sg13g2_decap_4
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_fill_2
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_720 VPWR VGND sg13g2_decap_8
XFILLER_0_263 VPWR VGND sg13g2_decap_8
XFILLER_1_797 VPWR VGND sg13g2_decap_8
XFILLER_49_779 VPWR VGND sg13g2_fill_2
XFILLER_36_418 VPWR VGND sg13g2_fill_2
XFILLER_45_985 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_fill_2
XFILLER_32_646 VPWR VGND sg13g2_decap_4
XFILLER_32_668 VPWR VGND sg13g2_decap_8
XFILLER_32_679 VPWR VGND sg13g2_fill_2
X_2740_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\] _0747_ _0506_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_178 VPWR VGND sg13g2_fill_2
XFILLER_9_875 VPWR VGND sg13g2_decap_8
XFILLER_12_392 VPWR VGND sg13g2_fill_2
X_2671_ _0734_ _0717_ _0731_ VPWR VGND sg13g2_nand2_2
X_4410_ net605 _2087_ _2101_ VPWR VGND sg13g2_and2_1
X_4341_ _2037_ _2017_ _2036_ VPWR VGND sg13g2_xnor2_1
X_4272_ _1977_ _1973_ _1976_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_3223_ net747 _0969_ _0970_ _0353_ VPWR VGND sg13g2_nor3_1
XFILLER_39_267 VPWR VGND sg13g2_fill_2
XFILLER_39_245 VPWR VGND sg13g2_decap_4
X_3154_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0923_ _0926_ VPWR VGND
+ sg13g2_nor2_1
X_3085_ _0875_ _0873_ _0874_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_123 VPWR VGND sg13g2_fill_1
XFILLER_11_819 VPWR VGND sg13g2_fill_2
X_3987_ _1713_ _1240_ _1711_ VPWR VGND sg13g2_nand2_1
XFILLER_23_679 VPWR VGND sg13g2_decap_4
XFILLER_10_329 VPWR VGND sg13g2_decap_8
X_2938_ videogen.fancy_shader.video_x\[3\] _0795_ _0796_ VPWR VGND sg13g2_and2_1
XFILLER_22_189 VPWR VGND sg13g2_decap_4
X_2869_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[2\] net762 _0778_ _0399_
+ VPWR VGND sg13g2_mux2_1
X_4608_ net691 net743 _0161_ VPWR VGND sg13g2_nor2_1
X_4539_ net680 net726 _0092_ VPWR VGND sg13g2_nor2_1
XFILLER_46_749 VPWR VGND sg13g2_fill_2
XFILLER_18_418 VPWR VGND sg13g2_decap_4
X_4843__311 VPWR VGND net311 sg13g2_tiehi
XFILLER_26_75 VPWR VGND sg13g2_decap_8
XFILLER_27_996 VPWR VGND sg13g2_decap_8
XFILLER_42_944 VPWR VGND sg13g2_decap_8
XFILLER_13_156 VPWR VGND sg13g2_fill_2
XFILLER_42_41 VPWR VGND sg13g2_fill_1
XFILLER_6_812 VPWR VGND sg13g2_decap_8
XFILLER_5_322 VPWR VGND sg13g2_decap_8
XFILLER_6_867 VPWR VGND sg13g2_fill_2
XFILLER_6_856 VPWR VGND sg13g2_decap_8
XFILLER_5_366 VPWR VGND sg13g2_decap_4
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_36_226 VPWR VGND sg13g2_decap_4
XFILLER_18_952 VPWR VGND sg13g2_decap_8
X_3910_ _1093_ _1632_ _1636_ VPWR VGND sg13g2_and2_1
X_4890_ net216 VGND VPWR _0441_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\]
+ _0098_ sg13g2_dfrbpq_1
XFILLER_32_410 VPWR VGND sg13g2_decap_8
X_3841_ VGND VPWR _1570_ net563 videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\]
+ sg13g2_or2_1
X_3772_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\] net564 _1502_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_34_1021 VPWR VGND sg13g2_decap_8
X_2723_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\] net769 _0744_ _0520_
+ VPWR VGND sg13g2_mux2_1
X_5511_ net600 net12 VPWR VGND sg13g2_buf_1
X_2654_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\] _0729_ _0574_
+ VPWR VGND sg13g2_mux2_1
X_2585_ _0689_ _0699_ _0700_ VPWR VGND sg13g2_nor2_2
X_4324_ net569 _2020_ _0619_ VPWR VGND sg13g2_nor2_1
X_4255_ VGND VPWR _1961_ _1960_ _0889_ sg13g2_or2_1
XFILLER_41_1014 VPWR VGND sg13g2_decap_8
X_3206_ videogen.fancy_shader.n646\[1\] _0957_ _0960_ VPWR VGND sg13g2_and2_1
X_4186_ VGND VPWR _0380_ _1905_ _0381_ sg13g2_or2_1
XFILLER_28_716 VPWR VGND sg13g2_decap_8
X_3137_ net748 _0912_ _0317_ VPWR VGND sg13g2_nor2_1
XFILLER_27_226 VPWR VGND sg13g2_decap_8
XFILLER_28_727 VPWR VGND sg13g2_fill_1
XFILLER_27_259 VPWR VGND sg13g2_decap_8
XFILLER_24_911 VPWR VGND sg13g2_decap_8
X_3068_ tmds_red.n114 tmds_red.n132 _0858_ VPWR VGND sg13g2_nor2_1
XFILLER_24_988 VPWR VGND sg13g2_decap_8
XFILLER_23_498 VPWR VGND sg13g2_fill_2
XFILLER_10_126 VPWR VGND sg13g2_fill_2
XFILLER_12_66 VPWR VGND sg13g2_fill_1
XFILLER_12_99 VPWR VGND sg13g2_decap_4
XFILLER_3_848 VPWR VGND sg13g2_decap_4
Xfanout651 net652 net651 VPWR VGND sg13g2_buf_8
Xfanout640 net642 net640 VPWR VGND sg13g2_buf_8
X_4810__354 VPWR VGND net354 sg13g2_tiehi
Xfanout662 net663 net662 VPWR VGND sg13g2_buf_1
Xfanout684 net693 net684 VPWR VGND sg13g2_buf_8
Xfanout673 net694 net673 VPWR VGND sg13g2_buf_8
Xfanout695 net696 net695 VPWR VGND sg13g2_buf_8
XFILLER_37_52 VPWR VGND sg13g2_fill_1
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_30_958 VPWR VGND sg13g2_decap_8
XFILLER_10_660 VPWR VGND sg13g2_decap_4
XFILLER_10_682 VPWR VGND sg13g2_decap_4
XFILLER_5_141 VPWR VGND sg13g2_fill_1
XFILLER_2_881 VPWR VGND sg13g2_decap_8
X_4040_ _1728_ _1749_ _1763_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_373 VPWR VGND sg13g2_decap_8
XFILLER_37_524 VPWR VGND sg13g2_decap_8
XFILLER_37_568 VPWR VGND sg13g2_fill_2
X_4942_ net61 VGND VPWR _0489_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\]
+ _0146_ sg13g2_dfrbpq_1
X_4873_ net249 VGND VPWR _0424_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\]
+ _0081_ sg13g2_dfrbpq_1
XFILLER_21_936 VPWR VGND sg13g2_decap_8
X_3824_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\] net579 _1553_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_446 VPWR VGND sg13g2_fill_2
X_3755_ net592 _1479_ _1484_ _1485_ VPWR VGND sg13g2_nor3_1
XFILLER_20_468 VPWR VGND sg13g2_fill_1
X_3686_ _1412_ _1413_ _1414_ _1415_ _1416_ VPWR VGND sg13g2_nor4_1
X_2706_ _0741_ _0706_ _0715_ VPWR VGND sg13g2_nand2_2
X_2637_ _0714_ _0723_ _0724_ VPWR VGND sg13g2_nor2_2
XFILLER_0_807 VPWR VGND sg13g2_decap_8
X_2568_ _0636_ _0681_ _0683_ VPWR VGND sg13g2_and2_1
X_4307_ _2000_ _2007_ _0615_ VPWR VGND sg13g2_nor2b_1
X_4238_ _1945_ _1944_ _1942_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_502 VPWR VGND sg13g2_decap_8
XFILLER_28_524 VPWR VGND sg13g2_decap_8
X_4169_ _1892_ _1235_ _1891_ VPWR VGND sg13g2_nand2_1
XFILLER_43_505 VPWR VGND sg13g2_fill_2
X_4907__182 VPWR VGND net182 sg13g2_tiehi
XFILLER_36_590 VPWR VGND sg13g2_decap_4
XFILLER_12_925 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_23_295 VPWR VGND sg13g2_decap_4
XFILLER_23_76 VPWR VGND sg13g2_fill_2
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_2_122 VPWR VGND sg13g2_fill_1
XFILLER_3_656 VPWR VGND sg13g2_decap_8
XFILLER_2_199 VPWR VGND sg13g2_fill_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_46_376 VPWR VGND sg13g2_fill_2
XFILLER_14_262 VPWR VGND sg13g2_decap_4
XFILLER_15_796 VPWR VGND sg13g2_fill_2
XFILLER_42_593 VPWR VGND sg13g2_decap_8
XFILLER_7_940 VPWR VGND sg13g2_decap_8
X_3540_ net619 VPWR _1270_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\]
+ net572 sg13g2_o21ai_1
XFILLER_11_991 VPWR VGND sg13g2_decap_8
XFILLER_6_472 VPWR VGND sg13g2_decap_4
X_3471_ _1200_ _1197_ _1066_ _1201_ VPWR VGND sg13g2_a21o_1
X_5072_ net146 VGND VPWR _0619_ tmds_green.dc_balancing_reg\[1\] net648 sg13g2_dfrbpq_2
X_4023_ _1735_ _1736_ _1739_ _1742_ _1746_ VPWR VGND sg13g2_nor4_1
XFILLER_49_181 VPWR VGND sg13g2_fill_2
XFILLER_37_354 VPWR VGND sg13g2_decap_8
XFILLER_25_516 VPWR VGND sg13g2_decap_4
XFILLER_37_398 VPWR VGND sg13g2_fill_1
XFILLER_25_549 VPWR VGND sg13g2_decap_4
X_4925_ net124 VGND VPWR _0476_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\]
+ _0133_ sg13g2_dfrbpq_1
X_4856_ net286 VGND VPWR _0407_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\]
+ _0064_ sg13g2_dfrbpq_1
XFILLER_20_232 VPWR VGND sg13g2_fill_1
XFILLER_21_766 VPWR VGND sg13g2_fill_1
X_3807_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\] net564 _1537_ VPWR
+ VGND sg13g2_nor2_1
X_4787_ net400 VGND VPWR _0338_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\]
+ _0038_ sg13g2_dfrbpq_1
X_3738_ net615 VPWR _1468_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\]
+ net551 sg13g2_o21ai_1
XFILLER_4_409 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_25 VPWR VGND uio_oe[4] sg13g2_tielo
X_3669_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1398_ _1399_ VPWR VGND
+ sg13g2_nor2_1
XFILLER_0_604 VPWR VGND sg13g2_decap_8
XFILLER_29_855 VPWR VGND sg13g2_fill_2
XFILLER_16_538 VPWR VGND sg13g2_fill_1
XFILLER_24_560 VPWR VGND sg13g2_decap_8
XFILLER_24_571 VPWR VGND sg13g2_fill_1
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_715 VPWR VGND sg13g2_decap_8
XFILLER_11_265 VPWR VGND sg13g2_fill_2
XFILLER_7_269 VPWR VGND sg13g2_fill_1
XFILLER_7_258 VPWR VGND sg13g2_fill_1
XFILLER_4_943 VPWR VGND sg13g2_decap_8
XFILLER_3_453 VPWR VGND sg13g2_decap_8
XFILLER_47_663 VPWR VGND sg13g2_decap_8
XFILLER_47_652 VPWR VGND sg13g2_fill_2
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_19_343 VPWR VGND sg13g2_decap_8
XFILLER_46_195 VPWR VGND sg13g2_fill_1
XFILLER_34_335 VPWR VGND sg13g2_fill_1
X_2971_ VPWR _0819_ _0818_ VGND sg13g2_inv_1
X_4710_ net653 net704 _0261_ VPWR VGND sg13g2_nor2_1
X_4641_ net661 net712 _0194_ VPWR VGND sg13g2_nor2_1
XFILLER_30_585 VPWR VGND sg13g2_decap_8
X_4572_ net685 net736 _0125_ VPWR VGND sg13g2_nor2_1
XFILLER_7_781 VPWR VGND sg13g2_decap_8
X_3523_ _1253_ net624 net626 VPWR VGND sg13g2_nand2b_1
X_3454_ _1147_ _1156_ _1183_ _1184_ VPWR VGND sg13g2_or3_1
X_3385_ _1088_ net542 _1115_ VPWR VGND sg13g2_nor2_1
X_5124_ net798 VGND VPWR serialize.n427\[8\] serialize.n411\[6\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5055_ net377 VGND VPWR _0602_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\]
+ _0250_ sg13g2_dfrbpq_1
X_4006_ _1039_ _1068_ _1725_ _1729_ VPWR VGND sg13g2_nor3_2
XFILLER_25_335 VPWR VGND sg13g2_fill_2
X_4908_ net180 VGND VPWR _0459_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\]
+ _0116_ sg13g2_dfrbpq_1
Xclkbuf_3_4__f_clk_regs clknet_0_clk_regs clknet_3_4__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_21_574 VPWR VGND sg13g2_decap_8
X_4839_ net319 VGND VPWR _0390_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\]
+ _0047_ sg13g2_dfrbpq_1
XFILLER_21_596 VPWR VGND sg13g2_decap_8
XFILLER_4_228 VPWR VGND sg13g2_decap_4
XFILLER_1_902 VPWR VGND sg13g2_decap_8
XFILLER_20_55 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_1_979 VPWR VGND sg13g2_decap_8
XFILLER_49_939 VPWR VGND sg13g2_decap_8
Xhold31 serialize.n417\[3\] VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold20 serialize.n414\[0\] VPWR VGND net425 sg13g2_dlygate4sd3_1
XFILLER_0_478 VPWR VGND sg13g2_fill_1
XFILLER_29_31 VPWR VGND sg13g2_decap_8
XFILLER_29_64 VPWR VGND sg13g2_decap_8
XFILLER_29_663 VPWR VGND sg13g2_fill_2
X_4881__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_28_151 VPWR VGND sg13g2_fill_1
XFILLER_28_162 VPWR VGND sg13g2_decap_4
XFILLER_45_63 VPWR VGND sg13g2_decap_4
XFILLER_45_52 VPWR VGND sg13g2_decap_8
XFILLER_43_143 VPWR VGND sg13g2_fill_2
XFILLER_31_305 VPWR VGND sg13g2_fill_1
XFILLER_39_416 VPWR VGND sg13g2_fill_1
X_3170_ net621 _0935_ _0937_ VPWR VGND sg13g2_nor2_1
XFILLER_39_427 VPWR VGND sg13g2_fill_2
XFILLER_48_972 VPWR VGND sg13g2_decap_8
XFILLER_35_633 VPWR VGND sg13g2_decap_4
XFILLER_47_493 VPWR VGND sg13g2_fill_1
XFILLER_22_316 VPWR VGND sg13g2_fill_1
XFILLER_15_390 VPWR VGND sg13g2_decap_8
X_2954_ VGND VPWR _0794_ _0811_ _0002_ _0371_ sg13g2_a21oi_1
X_2885_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\] net772 _0781_ _0343_
+ VPWR VGND sg13g2_mux2_1
X_4624_ net688 net740 _0177_ VPWR VGND sg13g2_nor2_1
X_4555_ net682 net733 _0108_ VPWR VGND sg13g2_nor2_1
X_3506_ _1236_ _1219_ _1233_ VPWR VGND sg13g2_xnor2_1
X_4486_ net685 net736 _0039_ VPWR VGND sg13g2_nor2_1
X_3437_ _1148_ _1155_ _1167_ VPWR VGND sg13g2_nor2_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_3368_ _1098_ videogen.fancy_shader.video_y\[9\] videogen.fancy_shader.n646\[9\]
+ VPWR VGND sg13g2_xnor2_1
X_5107_ net796 VGND VPWR serialize.n429\[4\] serialize.n417\[2\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_39_972 VPWR VGND sg13g2_decap_8
X_3299_ net611 videogen.fancy_shader.video_y\[3\] _1029_ VPWR VGND sg13g2_xor2_1
X_5038_ net236 VGND VPWR _0585_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\]
+ _0233_ sg13g2_dfrbpq_1
XFILLER_38_471 VPWR VGND sg13g2_decap_8
XFILLER_14_828 VPWR VGND sg13g2_fill_1
XFILLER_26_677 VPWR VGND sg13g2_decap_8
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_21_371 VPWR VGND sg13g2_decap_8
XFILLER_21_382 VPWR VGND sg13g2_fill_1
XFILLER_31_21 VPWR VGND sg13g2_fill_1
XFILLER_31_32 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
Xoutput8 net8 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_776 VPWR VGND sg13g2_decap_8
XFILLER_49_758 VPWR VGND sg13g2_fill_2
XFILLER_17_622 VPWR VGND sg13g2_decap_8
XFILLER_45_964 VPWR VGND sg13g2_decap_8
XFILLER_17_644 VPWR VGND sg13g2_fill_2
XFILLER_32_625 VPWR VGND sg13g2_decap_8
XFILLER_9_821 VPWR VGND sg13g2_decap_8
X_2670_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\] _0733_ _0562_
+ VPWR VGND sg13g2_mux2_1
X_4340_ _2034_ _2035_ _2036_ VPWR VGND sg13g2_nor2b_1
X_4271_ _1976_ tmds_red.dc_balancing_reg\[4\] _1975_ VPWR VGND sg13g2_xnor2_1
X_3222_ videogen.fancy_shader.n646\[7\] _0968_ _0970_ VPWR VGND sg13g2_and2_1
X_3153_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0923_ _0925_ VPWR VGND
+ sg13g2_and2_1
X_3084_ _0864_ VPWR _0874_ VGND net548 _0863_ sg13g2_o21ai_1
XFILLER_36_953 VPWR VGND sg13g2_decap_4
XFILLER_35_452 VPWR VGND sg13g2_fill_1
XFILLER_35_463 VPWR VGND sg13g2_fill_2
XFILLER_23_625 VPWR VGND sg13g2_decap_8
XFILLER_10_308 VPWR VGND sg13g2_decap_8
X_3986_ VGND VPWR _1702_ _1704_ _1712_ _1708_ sg13g2_a21oi_1
X_2937_ _0795_ videogen.fancy_shader.video_x\[2\] videogen.fancy_shader.video_x\[1\]
+ net630 VPWR VGND sg13g2_and3_2
X_4607_ net691 net743 _0160_ VPWR VGND sg13g2_nor2_1
X_2868_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\] net752 _0778_ _0400_
+ VPWR VGND sg13g2_mux2_1
X_2799_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\] _0760_ _0451_
+ VPWR VGND sg13g2_mux2_1
X_4538_ net679 net730 _0091_ VPWR VGND sg13g2_nor2_1
Xfanout800 net802 net800 VPWR VGND sg13g2_buf_8
X_4469_ net661 net712 _0022_ VPWR VGND sg13g2_nor2_1
XFILLER_42_923 VPWR VGND sg13g2_decap_8
XFILLER_27_975 VPWR VGND sg13g2_decap_8
XFILLER_26_485 VPWR VGND sg13g2_decap_8
XFILLER_9_128 VPWR VGND sg13g2_decap_4
XFILLER_42_86 VPWR VGND sg13g2_decap_8
X_4917__162 VPWR VGND net162 sg13g2_tiehi
X_4733__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_3_36 VPWR VGND sg13g2_fill_1
XFILLER_49_511 VPWR VGND sg13g2_decap_8
XFILLER_37_706 VPWR VGND sg13g2_decap_8
XFILLER_3_1009 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_36_205 VPWR VGND sg13g2_decap_8
XFILLER_18_931 VPWR VGND sg13g2_decap_8
XFILLER_33_901 VPWR VGND sg13g2_decap_8
X_3840_ VGND VPWR _1569_ net553 videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\]
+ sg13g2_or2_1
XFILLER_34_1000 VPWR VGND sg13g2_decap_8
X_3771_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\] net577 _1501_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_13_680 VPWR VGND sg13g2_decap_4
X_2722_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\] net759 _0744_ _0521_
+ VPWR VGND sg13g2_mux2_1
X_5510_ videogen.mem_row net11 VPWR VGND sg13g2_buf_8
X_2653_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\] _0729_ _0575_
+ VPWR VGND sg13g2_mux2_1
X_2584_ _0699_ _0696_ _0697_ VPWR VGND sg13g2_nand2_2
X_4323_ _2020_ _0642_ _2019_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_890 VPWR VGND sg13g2_decap_8
X_4254_ _1940_ _1959_ _1960_ VPWR VGND sg13g2_nor2_1
X_3205_ videogen.fancy_shader.n646\[1\] _0957_ _0959_ VPWR VGND sg13g2_nor2_1
X_4185_ VGND VPWR _0379_ _1906_ _0381_ sg13g2_or2_1
X_3136_ _0662_ _0663_ _0814_ _0911_ _0912_ VPWR VGND sg13g2_nor4_1
X_3067_ _0857_ tmds_red.n114 tmds_red.n132 VPWR VGND sg13g2_nand2_1
XFILLER_23_455 VPWR VGND sg13g2_decap_4
XFILLER_24_967 VPWR VGND sg13g2_decap_8
X_4899__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_23_488 VPWR VGND sg13g2_decap_4
X_3969_ _1692_ _1693_ _1690_ _1695_ VPWR VGND sg13g2_nand3_1
XFILLER_12_23 VPWR VGND sg13g2_decap_8
X_4953__395 VPWR VGND net395 sg13g2_tiehi
XFILLER_2_348 VPWR VGND sg13g2_fill_1
XFILLER_2_359 VPWR VGND sg13g2_decap_8
Xfanout641 net642 net641 VPWR VGND sg13g2_buf_8
Xfanout630 videogen.fancy_shader.video_x\[0\] net630 VPWR VGND sg13g2_buf_8
Xfanout652 net656 net652 VPWR VGND sg13g2_buf_8
Xfanout674 net678 net674 VPWR VGND sg13g2_buf_8
Xfanout663 net673 net663 VPWR VGND sg13g2_buf_8
Xfanout685 net693 net685 VPWR VGND sg13g2_buf_8
Xfanout696 net430 net696 VPWR VGND sg13g2_buf_8
XFILLER_46_547 VPWR VGND sg13g2_fill_1
XFILLER_46_536 VPWR VGND sg13g2_decap_8
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_33_219 VPWR VGND sg13g2_fill_1
XFILLER_41_274 VPWR VGND sg13g2_fill_2
XFILLER_41_252 VPWR VGND sg13g2_decap_4
XFILLER_30_937 VPWR VGND sg13g2_decap_8
XFILLER_6_687 VPWR VGND sg13g2_fill_2
XFILLER_6_676 VPWR VGND sg13g2_fill_1
XFILLER_45_7 VPWR VGND sg13g2_fill_2
XFILLER_2_860 VPWR VGND sg13g2_decap_8
X_4711__253 VPWR VGND net253 sg13g2_tiehi
XFILLER_49_352 VPWR VGND sg13g2_decap_8
X_4941_ net65 VGND VPWR _0488_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\]
+ _0145_ sg13g2_dfrbpq_1
X_4872_ net251 VGND VPWR _0423_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\]
+ _0080_ sg13g2_dfrbpq_1
X_3823_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\] net565 _1552_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_21_915 VPWR VGND sg13g2_decap_8
XFILLER_33_786 VPWR VGND sg13g2_fill_2
X_3754_ _1480_ _1481_ _1482_ _1483_ _1484_ VPWR VGND sg13g2_nor4_1
X_3685_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[1\] net582 _1415_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_492 VPWR VGND sg13g2_fill_2
X_2705_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\] _0740_ _0534_
+ VPWR VGND sg13g2_mux2_1
X_2636_ net592 _0693_ _0709_ _0723_ VPWR VGND sg13g2_or3_1
X_2567_ _0682_ net612 _0676_ VPWR VGND sg13g2_xnor2_1
X_4306_ _2005_ _2006_ _2001_ _2007_ VPWR VGND sg13g2_mux2_1
X_4237_ _0855_ _1929_ _1944_ VPWR VGND sg13g2_nor2_1
X_4168_ _1878_ VPWR _1891_ VGND _1856_ _1870_ sg13g2_o21ai_1
X_4099_ _1818_ _1820_ _1813_ _1822_ VPWR VGND sg13g2_nand3_1
X_3119_ _0796_ _0901_ _0306_ VPWR VGND sg13g2_nor2_1
XFILLER_15_219 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_8_919 VPWR VGND sg13g2_decap_8
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_fill_2
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_19_558 VPWR VGND sg13g2_fill_1
XFILLER_15_753 VPWR VGND sg13g2_decap_4
X_4995__215 VPWR VGND net215 sg13g2_tiehi
XFILLER_9_57 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_31_1025 VPWR VGND sg13g2_decap_4
XFILLER_7_996 VPWR VGND sg13g2_decap_8
X_3470_ _1190_ VPWR _1200_ VGND _1198_ _1199_ sg13g2_o21ai_1
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_5028__318 VPWR VGND net318 sg13g2_tiehi
X_5071_ net161 VGND VPWR _0618_ blue_tmds_par\[9\] net641 sg13g2_dfrbpq_1
XFILLER_38_812 VPWR VGND sg13g2_decap_4
X_4022_ VPWR VGND _1741_ _1736_ _1739_ _1733_ _1745_ _1734_ sg13g2_a221oi_1
XFILLER_49_160 VPWR VGND sg13g2_decap_8
XFILLER_38_856 VPWR VGND sg13g2_fill_2
XFILLER_38_878 VPWR VGND sg13g2_decap_4
Xclkbuf_3_3__f_clk_regs clknet_0_clk_regs clknet_3_3__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_40_509 VPWR VGND sg13g2_decap_4
X_4924_ net128 VGND VPWR _0475_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\]
+ _0132_ sg13g2_dfrbpq_1
X_4855_ net288 VGND VPWR _0406_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\]
+ _0063_ sg13g2_dfrbpq_1
XFILLER_20_200 VPWR VGND sg13g2_decap_4
X_4786_ net404 VGND VPWR _0337_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\]
+ net634 sg13g2_dfrbpq_1
X_3806_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\] net586 _1536_ VPWR
+ VGND sg13g2_nor2_1
X_3737_ _1463_ _1464_ _1465_ _1466_ _1467_ VPWR VGND sg13g2_nor4_1
Xheichips25_bagel_26 VPWR VGND uio_oe[5] sg13g2_tielo
X_3668_ net612 _1386_ _1397_ _1398_ VPWR VGND sg13g2_nor3_1
X_3599_ _1325_ _1326_ _1327_ _1328_ _1329_ VPWR VGND sg13g2_nor4_1
X_2619_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\] _0716_ _0596_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_627 VPWR VGND sg13g2_fill_1
XFILLER_0_649 VPWR VGND sg13g2_decap_8
XFILLER_18_22 VPWR VGND sg13g2_fill_2
XFILLER_18_77 VPWR VGND sg13g2_fill_1
XFILLER_44_837 VPWR VGND sg13g2_decap_8
XFILLER_28_388 VPWR VGND sg13g2_fill_2
XFILLER_12_712 VPWR VGND sg13g2_decap_8
XFILLER_12_723 VPWR VGND sg13g2_fill_1
XFILLER_4_922 VPWR VGND sg13g2_decap_8
XFILLER_4_999 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_4
XFILLER_3_498 VPWR VGND sg13g2_fill_1
X_4851__296 VPWR VGND net296 sg13g2_tiehi
XFILLER_19_300 VPWR VGND sg13g2_decap_4
XFILLER_46_185 VPWR VGND sg13g2_fill_2
XFILLER_19_399 VPWR VGND sg13g2_decap_8
XFILLER_34_325 VPWR VGND sg13g2_fill_2
X_2970_ _0665_ _0817_ _0818_ VPWR VGND sg13g2_nor2_2
XFILLER_30_520 VPWR VGND sg13g2_fill_2
X_4640_ net666 net718 _0193_ VPWR VGND sg13g2_nor2_1
X_4571_ net677 net729 _0124_ VPWR VGND sg13g2_nor2_1
X_3522_ net619 VPWR _1252_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\]
+ net583 sg13g2_o21ai_1
X_3453_ VPWR VGND _1168_ _1158_ _1166_ _1019_ _1183_ _1020_ sg13g2_a221oi_1
X_3384_ VPWR _1114_ _1113_ VGND sg13g2_inv_1
XFILLER_34_0 VPWR VGND sg13g2_decap_4
X_5123_ net798 VGND VPWR serialize.n427\[7\] serialize.n411\[5\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5054_ net39 VGND VPWR _0601_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\]
+ _0249_ sg13g2_dfrbpq_1
X_5080__353 VPWR VGND net353 sg13g2_tiehi
XFILLER_37_130 VPWR VGND sg13g2_decap_4
X_4005_ _1728_ _1659_ _1726_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_815 VPWR VGND sg13g2_decap_8
XFILLER_25_358 VPWR VGND sg13g2_decap_4
XFILLER_40_317 VPWR VGND sg13g2_fill_1
X_4907_ net182 VGND VPWR _0458_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\]
+ _0115_ sg13g2_dfrbpq_1
XFILLER_33_391 VPWR VGND sg13g2_fill_2
X_4838_ net321 VGND VPWR _0389_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\]
+ _0046_ sg13g2_dfrbpq_1
XFILLER_21_553 VPWR VGND sg13g2_decap_8
XFILLER_14_1020 VPWR VGND sg13g2_decap_8
X_4769_ net64 VGND VPWR _0320_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\]
+ net631 sg13g2_dfrbpq_1
XFILLER_1_958 VPWR VGND sg13g2_decap_8
XFILLER_49_918 VPWR VGND sg13g2_decap_8
Xhold21 serialize.n417\[1\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold10 serialize.n420\[6\] VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold32 serialize.n411\[3\] VPWR VGND net437 sg13g2_dlygate4sd3_1
X_4985__258 VPWR VGND net258 sg13g2_tiehi
XFILLER_21_1013 VPWR VGND sg13g2_decap_8
XFILLER_28_141 VPWR VGND sg13g2_fill_1
XFILLER_16_314 VPWR VGND sg13g2_decap_4
XFILLER_29_675 VPWR VGND sg13g2_decap_4
XFILLER_44_645 VPWR VGND sg13g2_fill_2
XFILLER_43_133 VPWR VGND sg13g2_fill_2
XFILLER_44_678 VPWR VGND sg13g2_fill_2
XFILLER_43_177 VPWR VGND sg13g2_fill_2
XFILLER_25_892 VPWR VGND sg13g2_decap_8
XFILLER_4_763 VPWR VGND sg13g2_fill_2
XFILLER_48_951 VPWR VGND sg13g2_decap_8
X_4743__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_35_656 VPWR VGND sg13g2_fill_2
X_2953_ _0807_ _0808_ net793 _0811_ VPWR VGND _0809_ sg13g2_nand4_1
XFILLER_16_881 VPWR VGND sg13g2_decap_8
X_2884_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\] net762 _0781_ _0344_
+ VPWR VGND sg13g2_mux2_1
X_4623_ net689 net742 _0176_ VPWR VGND sg13g2_nor2_1
X_4554_ net682 net733 _0107_ VPWR VGND sg13g2_nor2_1
X_3505_ net630 videogen.fancy_shader.video_y\[0\] _1235_ VPWR VGND sg13g2_xor2_1
X_4485_ net686 net737 _0038_ VPWR VGND sg13g2_nor2_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_3436_ _1162_ _1163_ _1160_ _1166_ VPWR VGND sg13g2_nand3_1
X_3367_ _1089_ VPWR _1097_ VGND _1094_ _1095_ sg13g2_o21ai_1
X_5106_ net800 VGND VPWR serialize.n429\[3\] serialize.n417\[1\] clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5037_ net244 VGND VPWR _0584_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\]
+ _0232_ sg13g2_dfrbpq_1
X_3298_ videogen.fancy_shader.video_y\[3\] net611 _1028_ VPWR VGND sg13g2_nor2_1
XFILLER_13_306 VPWR VGND sg13g2_decap_4
XFILLER_25_155 VPWR VGND sg13g2_fill_2
XFILLER_25_199 VPWR VGND sg13g2_fill_2
XFILLER_5_516 VPWR VGND sg13g2_fill_2
Xoutput9 net9 uio_out[3] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_755 VPWR VGND sg13g2_decap_8
XFILLER_49_737 VPWR VGND sg13g2_decap_8
XFILLER_45_943 VPWR VGND sg13g2_decap_8
XFILLER_44_431 VPWR VGND sg13g2_decap_4
XFILLER_17_689 VPWR VGND sg13g2_fill_1
XFILLER_13_851 VPWR VGND sg13g2_fill_1
XFILLER_31_158 VPWR VGND sg13g2_decap_8
XFILLER_13_884 VPWR VGND sg13g2_decap_4
XFILLER_9_855 VPWR VGND sg13g2_decap_4
X_4270_ VGND VPWR tmds_red.dc_balancing_reg\[3\] _1954_ _1975_ _1974_ sg13g2_a21oi_1
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
X_3221_ videogen.fancy_shader.n646\[7\] _0968_ _0969_ VPWR VGND sg13g2_nor2_1
X_3152_ _0919_ _0923_ _0924_ _0320_ VPWR VGND sg13g2_nor3_1
XFILLER_39_269 VPWR VGND sg13g2_fill_1
X_3083_ _0869_ _0861_ _0872_ _0873_ VPWR VGND sg13g2_a21o_1
XFILLER_36_921 VPWR VGND sg13g2_decap_8
XFILLER_48_792 VPWR VGND sg13g2_decap_4
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_23_604 VPWR VGND sg13g2_decap_8
X_3985_ _1694_ _1697_ _1690_ _1711_ VPWR VGND sg13g2_mux2_1
XFILLER_22_158 VPWR VGND sg13g2_decap_8
X_2936_ _0794_ _0793_ VPWR VGND sg13g2_inv_2
X_2867_ _0723_ _0772_ _0778_ VPWR VGND sg13g2_nor2_2
X_4606_ net691 net743 _0159_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
X_2798_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[3\] _0760_ _0452_
+ VPWR VGND sg13g2_mux2_1
X_4537_ net679 net726 _0090_ VPWR VGND sg13g2_nor2_1
X_4468_ net674 net726 _0021_ VPWR VGND sg13g2_nor2_1
Xfanout801 net802 net801 VPWR VGND sg13g2_buf_8
X_3419_ VPWR VGND _1143_ _1134_ _1141_ _1053_ _1149_ _1054_ sg13g2_a221oi_1
X_4399_ VPWR _2090_ _2089_ VGND sg13g2_inv_1
XFILLER_39_781 VPWR VGND sg13g2_decap_4
XFILLER_27_954 VPWR VGND sg13g2_decap_8
XFILLER_42_902 VPWR VGND sg13g2_decap_8
XFILLER_26_44 VPWR VGND sg13g2_decap_8
XFILLER_26_55 VPWR VGND sg13g2_fill_2
XFILLER_41_423 VPWR VGND sg13g2_fill_2
XFILLER_41_412 VPWR VGND sg13g2_decap_8
XFILLER_42_979 VPWR VGND sg13g2_decap_8
XFILLER_41_456 VPWR VGND sg13g2_decap_8
XFILLER_13_136 VPWR VGND sg13g2_fill_2
XFILLER_10_821 VPWR VGND sg13g2_decap_4
XFILLER_10_854 VPWR VGND sg13g2_fill_2
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_29_280 VPWR VGND sg13g2_decap_4
XFILLER_29_291 VPWR VGND sg13g2_fill_2
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_44_261 VPWR VGND sg13g2_fill_1
XFILLER_32_423 VPWR VGND sg13g2_fill_1
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_fill_2
XFILLER_33_979 VPWR VGND sg13g2_decap_8
X_3770_ net617 VPWR _1500_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\]
+ net586 sg13g2_o21ai_1
X_2721_ _0707_ _0723_ _0744_ VPWR VGND sg13g2_nor2_2
X_2652_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\] _0729_ _0576_
+ VPWR VGND sg13g2_mux2_1
X_2583_ _0696_ _0697_ _0698_ VPWR VGND sg13g2_and2_1
X_4322_ _2017_ _2018_ _2019_ VPWR VGND sg13g2_and2_1
X_4253_ _1957_ _1953_ _1959_ VPWR VGND sg13g2_xor2_1
X_3204_ _0957_ _0958_ _0346_ VPWR VGND sg13g2_nor2b_1
X_4184_ _1352_ _1550_ _1720_ _1906_ VPWR VGND sg13g2_nor3_1
X_3135_ _0911_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\]
+ VPWR VGND sg13g2_nand2b_1
X_3066_ tmds_red.dc_balancing_reg\[1\] tmds_red.dc_balancing_reg\[0\] tmds_red.dc_balancing_reg\[3\]
+ tmds_red.dc_balancing_reg\[2\] _0856_ VPWR VGND sg13g2_nor4_1
XFILLER_24_946 VPWR VGND sg13g2_decap_8
XFILLER_35_250 VPWR VGND sg13g2_fill_1
X_3968_ _1694_ _1692_ _1693_ VPWR VGND sg13g2_nand2_1
X_2919_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\] net763 _0788_ _0285_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_990 VPWR VGND sg13g2_decap_8
X_3899_ _1625_ _1175_ _1624_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_46 VPWR VGND sg13g2_fill_1
XFILLER_12_57 VPWR VGND sg13g2_decap_8
XFILLER_12_79 VPWR VGND sg13g2_fill_1
Xfanout642 net643 net642 VPWR VGND sg13g2_buf_8
Xfanout631 net632 net631 VPWR VGND sg13g2_buf_8
Xfanout620 net623 net620 VPWR VGND sg13g2_buf_8
Xfanout664 net667 net664 VPWR VGND sg13g2_buf_8
Xfanout675 net678 net675 VPWR VGND sg13g2_buf_8
Xfanout653 net655 net653 VPWR VGND sg13g2_buf_8
Xfanout697 net701 net697 VPWR VGND sg13g2_buf_8
Xfanout686 net687 net686 VPWR VGND sg13g2_buf_8
XFILLER_2_1021 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_fill_2
XFILLER_37_87 VPWR VGND sg13g2_fill_1
XFILLER_27_740 VPWR VGND sg13g2_fill_2
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_42_743 VPWR VGND sg13g2_fill_2
XFILLER_26_294 VPWR VGND sg13g2_fill_2
X_4878__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_14_467 VPWR VGND sg13g2_decap_8
XFILLER_14_478 VPWR VGND sg13g2_fill_1
XFILLER_30_916 VPWR VGND sg13g2_decap_8
XFILLER_41_286 VPWR VGND sg13g2_fill_2
X_4767__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_23_990 VPWR VGND sg13g2_decap_8
X_4782__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_6_633 VPWR VGND sg13g2_fill_1
XFILLER_5_110 VPWR VGND sg13g2_fill_1
XFILLER_49_331 VPWR VGND sg13g2_decap_8
Xclkbuf_3_2__f_clk_regs clknet_0_clk_regs clknet_3_2__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_4940_ net70 VGND VPWR _0487_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\]
+ _0144_ sg13g2_dfrbpq_1
XFILLER_18_773 VPWR VGND sg13g2_fill_2
XFILLER_18_795 VPWR VGND sg13g2_fill_1
X_4861__276 VPWR VGND net276 sg13g2_tiehi
X_4871_ net257 VGND VPWR _0422_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\]
+ _0079_ sg13g2_dfrbpq_1
X_3822_ VPWR _0372_ _1551_ VGND sg13g2_inv_1
XFILLER_33_798 VPWR VGND sg13g2_decap_4
XFILLER_20_448 VPWR VGND sg13g2_fill_1
X_3753_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\] net582 _1483_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_459 VPWR VGND sg13g2_decap_8
X_3684_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\] net559 _1414_ VPWR
+ VGND sg13g2_nor2_1
X_2704_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\] _0740_ _0535_
+ VPWR VGND sg13g2_mux2_1
X_2635_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\] net784 _0722_ _0586_
+ VPWR VGND sg13g2_mux2_1
X_4305_ _0647_ _2002_ _2004_ _2006_ VPWR VGND sg13g2_or3_1
X_2566_ _0637_ _0676_ _0681_ VPWR VGND sg13g2_and2_1
X_4236_ _1929_ _1942_ _1943_ VPWR VGND sg13g2_nor2_1
X_4167_ _1883_ _1875_ _1890_ VPWR VGND sg13g2_xor2_1
X_3118_ net795 VPWR _0901_ VGND videogen.fancy_shader.video_x\[3\] _0795_ sg13g2_o21ai_1
X_4098_ VPWR _1821_ _1820_ VGND sg13g2_inv_1
X_3049_ _0642_ _0839_ _0840_ VPWR VGND sg13g2_and2_1
XFILLER_24_754 VPWR VGND sg13g2_fill_2
XFILLER_11_415 VPWR VGND sg13g2_fill_2
XFILLER_23_253 VPWR VGND sg13g2_fill_2
XFILLER_3_614 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_146 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_48_75 VPWR VGND sg13g2_decap_4
XFILLER_19_515 VPWR VGND sg13g2_decap_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_46_323 VPWR VGND sg13g2_decap_4
XFILLER_46_301 VPWR VGND sg13g2_decap_4
XFILLER_34_529 VPWR VGND sg13g2_decap_8
X_4921__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_42_573 VPWR VGND sg13g2_fill_2
XFILLER_15_798 VPWR VGND sg13g2_fill_1
XFILLER_31_1004 VPWR VGND sg13g2_decap_8
XFILLER_10_470 VPWR VGND sg13g2_fill_1
X_4891__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_7_975 VPWR VGND sg13g2_decap_8
X_4791__392 VPWR VGND net392 sg13g2_tiehi
X_5070_ net169 VGND VPWR _0617_ blue_tmds_par\[8\] net642 sg13g2_dfrbpq_1
X_4021_ VPWR _1744_ _1743_ VGND sg13g2_inv_1
XFILLER_49_183 VPWR VGND sg13g2_fill_1
XFILLER_25_507 VPWR VGND sg13g2_decap_4
X_4923_ net132 VGND VPWR _0474_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\]
+ _0131_ sg13g2_dfrbpq_1
X_4854_ net290 VGND VPWR _0405_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\]
+ _0062_ sg13g2_dfrbpq_1
X_4785_ net32 VGND VPWR _0336_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\]
+ net633 sg13g2_dfrbpq_2
XFILLER_21_757 VPWR VGND sg13g2_decap_8
X_3805_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\] net554 _1535_ VPWR
+ VGND sg13g2_nor2_1
X_3736_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\] net575 _1466_ VPWR
+ VGND sg13g2_nor2_1
X_3667_ net620 _1391_ _1396_ _1397_ VPWR VGND sg13g2_nor3_1
Xheichips25_bagel_27 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_3598_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\] net552 _1328_ VPWR
+ VGND sg13g2_nor2_1
X_2618_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\] _0716_ _0597_
+ VPWR VGND sg13g2_mux2_1
X_2549_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\] net608
+ net609 _0664_ VPWR VGND sg13g2_nor4_1
X_4219_ tmds_red.dc_balancing_reg\[0\] _0836_ _0501_ VPWR VGND sg13g2_and2_1
XFILLER_28_312 VPWR VGND sg13g2_decap_8
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_18_45 VPWR VGND sg13g2_decap_8
XFILLER_16_518 VPWR VGND sg13g2_decap_8
XFILLER_16_529 VPWR VGND sg13g2_decap_8
XFILLER_7_249 VPWR VGND sg13g2_decap_8
XFILLER_4_901 VPWR VGND sg13g2_decap_8
XFILLER_4_978 VPWR VGND sg13g2_decap_8
XFILLER_19_378 VPWR VGND sg13g2_decap_8
XFILLER_35_827 VPWR VGND sg13g2_decap_8
XFILLER_34_359 VPWR VGND sg13g2_fill_2
XFILLER_15_562 VPWR VGND sg13g2_decap_4
XFILLER_43_893 VPWR VGND sg13g2_decap_8
X_4570_ net684 net735 _0123_ VPWR VGND sg13g2_nor2_1
X_3521_ net797 net1 _1251_ VPWR VGND sg13g2_and2_1
XFILLER_6_293 VPWR VGND sg13g2_fill_2
X_3452_ _1172_ _1181_ _1171_ _1182_ VPWR VGND sg13g2_nand3_1
X_3383_ _1113_ _1088_ net542 VPWR VGND sg13g2_nand2_1
X_5122_ net798 VGND VPWR net420 serialize.n411\[4\] clknet_3_4__leaf_clk_regs sg13g2_dfrbpq_1
X_5053_ net55 VGND VPWR _0600_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\]
+ _0248_ sg13g2_dfrbpq_1
X_4004_ VPWR _1727_ _1726_ VGND sg13g2_inv_1
XFILLER_40_329 VPWR VGND sg13g2_decap_8
X_4906_ net184 VGND VPWR _0457_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\]
+ _0114_ sg13g2_dfrbpq_1
XFILLER_21_532 VPWR VGND sg13g2_fill_1
X_4837_ net322 VGND VPWR _0388_ red_tmds_par\[9\] net644 sg13g2_dfrbpq_1
X_4768_ net66 VGND VPWR _0319_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\]
+ net631 sg13g2_dfrbpq_2
X_4699_ net691 net743 _0252_ VPWR VGND sg13g2_nor2_1
X_3719_ _1449_ _1400_ _1448_ _0650_ videogen.test_lut_thingy.gol_counter_reg\[1\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_20_68 VPWR VGND sg13g2_decap_4
XFILLER_0_403 VPWR VGND sg13g2_decap_8
XFILLER_1_937 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_4
Xhold11 serialize.n431\[6\] VPWR VGND net416 sg13g2_dlygate4sd3_1
XFILLER_48_407 VPWR VGND sg13g2_fill_2
Xhold22 serialize.n414\[6\] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold33 serialize.n411\[0\] VPWR VGND net438 sg13g2_dlygate4sd3_1
XFILLER_29_99 VPWR VGND sg13g2_fill_2
XFILLER_29_665 VPWR VGND sg13g2_fill_1
XFILLER_16_304 VPWR VGND sg13g2_decap_4
XFILLER_45_32 VPWR VGND sg13g2_fill_2
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_45_87 VPWR VGND sg13g2_decap_8
XFILLER_25_871 VPWR VGND sg13g2_decap_8
XFILLER_40_830 VPWR VGND sg13g2_fill_1
XFILLER_24_370 VPWR VGND sg13g2_fill_1
X_5057__345 VPWR VGND net345 sg13g2_tiehi
XFILLER_8_503 VPWR VGND sg13g2_decap_4
XFILLER_6_59 VPWR VGND sg13g2_fill_2
XFILLER_4_786 VPWR VGND sg13g2_decap_8
XFILLER_6_1019 VPWR VGND sg13g2_decap_4
XFILLER_48_930 VPWR VGND sg13g2_decap_8
XFILLER_23_819 VPWR VGND sg13g2_decap_8
XFILLER_35_668 VPWR VGND sg13g2_decap_8
X_2952_ _0810_ net793 _0809_ VPWR VGND sg13g2_nand2_1
X_2883_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\] net752 _0781_ _0345_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_351 VPWR VGND sg13g2_decap_8
XFILLER_30_362 VPWR VGND sg13g2_fill_1
XFILLER_30_395 VPWR VGND sg13g2_decap_4
X_4622_ net688 net740 _0175_ VPWR VGND sg13g2_nor2_1
X_4553_ net682 net733 _0106_ VPWR VGND sg13g2_nor2_1
X_4484_ net670 net721 _0037_ VPWR VGND sg13g2_nor2_1
XFILLER_7_580 VPWR VGND sg13g2_decap_8
X_3504_ _1234_ net609 net630 VPWR VGND sg13g2_xnor2_1
X_3435_ _1165_ _1160_ _1162_ _1163_ VPWR VGND sg13g2_and3_1
X_3366_ net610 videogen.fancy_shader.video_y\[8\] _1096_ VPWR VGND sg13g2_xor2_1
X_5105_ net800 VGND VPWR serialize.n429\[2\] serialize.n417\[0\] clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3297_ _1027_ _1025_ _1026_ VPWR VGND sg13g2_xnor2_1
X_5036_ net252 VGND VPWR _0583_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\]
+ _0231_ sg13g2_dfrbpq_1
XFILLER_14_819 VPWR VGND sg13g2_decap_8
XFILLER_15_13 VPWR VGND sg13g2_fill_2
XFILLER_41_627 VPWR VGND sg13g2_fill_1
XFILLER_15_57 VPWR VGND sg13g2_decap_4
XFILLER_21_362 VPWR VGND sg13g2_decap_4
XFILLER_31_12 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_200 VPWR VGND sg13g2_fill_1
XFILLER_1_734 VPWR VGND sg13g2_decap_8
XFILLER_0_244 VPWR VGND sg13g2_fill_1
XFILLER_0_277 VPWR VGND sg13g2_decap_8
XFILLER_45_922 VPWR VGND sg13g2_decap_8
XFILLER_17_646 VPWR VGND sg13g2_fill_1
XFILLER_45_999 VPWR VGND sg13g2_decap_8
XFILLER_31_137 VPWR VGND sg13g2_decap_8
XFILLER_8_355 VPWR VGND sg13g2_fill_1
XFILLER_8_388 VPWR VGND sg13g2_fill_2
XFILLER_9_889 VPWR VGND sg13g2_fill_2
XFILLER_4_572 VPWR VGND sg13g2_decap_8
X_3220_ net748 _0967_ _0968_ _0352_ VPWR VGND sg13g2_nor3_1
X_3151_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0922_ _0924_ VPWR VGND
+ sg13g2_nor2_1
X_3082_ _0861_ _0871_ _0872_ VPWR VGND sg13g2_nor2_1
XFILLER_35_476 VPWR VGND sg13g2_decap_8
XFILLER_35_487 VPWR VGND sg13g2_fill_2
X_3984_ _1710_ _1708_ _1709_ VPWR VGND sg13g2_nand2_1
X_2935_ _0793_ net793 VPWR VGND videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ sg13g2_nand2b_2
X_2866_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\] net785 _0777_ _0401_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_181 VPWR VGND sg13g2_fill_1
XFILLER_31_693 VPWR VGND sg13g2_fill_2
X_4605_ net691 net743 _0158_ VPWR VGND sg13g2_nor2_1
X_2797_ _0760_ _0698_ _0751_ VPWR VGND sg13g2_nand2_2
X_4536_ net657 net709 _0089_ VPWR VGND sg13g2_nor2_1
X_4467_ net675 net727 _0020_ VPWR VGND sg13g2_nor2_1
Xfanout802 net803 net802 VPWR VGND sg13g2_buf_8
X_3418_ _1036_ _1134_ _1145_ _1146_ _1148_ VPWR VGND sg13g2_nor4_1
X_4398_ _2083_ VPWR _2089_ VGND _0645_ _2076_ sg13g2_o21ai_1
X_3349_ _1078_ VPWR _1079_ VGND videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.n646\[5\]
+ sg13g2_o21ai_1
X_5019_ net59 VGND VPWR _0566_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\]
+ _0214_ sg13g2_dfrbpq_1
XFILLER_27_933 VPWR VGND sg13g2_decap_8
XFILLER_38_292 VPWR VGND sg13g2_fill_2
X_4779__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_26_89 VPWR VGND sg13g2_decap_4
XFILLER_42_958 VPWR VGND sg13g2_decap_8
XFILLER_42_11 VPWR VGND sg13g2_fill_2
XFILLER_41_435 VPWR VGND sg13g2_decap_8
XFILLER_41_479 VPWR VGND sg13g2_decap_8
XFILLER_42_66 VPWR VGND sg13g2_fill_2
XFILLER_22_682 VPWR VGND sg13g2_fill_1
XFILLER_5_347 VPWR VGND sg13g2_fill_1
XFILLER_3_27 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
X_4998__203 VPWR VGND net203 sg13g2_tiehi
XFILLER_45_752 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk_regs clknet_0_clk_regs clknet_3_1__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_18_966 VPWR VGND sg13g2_decap_8
XFILLER_44_273 VPWR VGND sg13g2_decap_4
XFILLER_32_402 VPWR VGND sg13g2_decap_4
XFILLER_33_947 VPWR VGND sg13g2_fill_2
XFILLER_33_958 VPWR VGND sg13g2_decap_8
XFILLER_20_608 VPWR VGND sg13g2_decap_4
X_2720_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\] _0743_ _0522_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_631 VPWR VGND sg13g2_fill_2
XFILLER_12_181 VPWR VGND sg13g2_decap_8
X_2651_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\] _0729_ _0577_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_152 VPWR VGND sg13g2_decap_4
XFILLER_12_192 VPWR VGND sg13g2_fill_2
X_2582_ VGND VPWR _0649_ _0697_ net543 net626 sg13g2_a21oi_2
X_4321_ _2016_ _2015_ net602 _2018_ VPWR VGND sg13g2_a21o_1
X_4252_ _1953_ _1957_ _1958_ VPWR VGND sg13g2_nor2b_1
X_3203_ VGND VPWR _0635_ _0918_ _0958_ net751 sg13g2_a21oi_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_4183_ _1550_ _1901_ _1905_ VPWR VGND sg13g2_nor2_1
X_3134_ _0898_ _0910_ _0312_ VPWR VGND sg13g2_nor2_1
XFILLER_48_590 VPWR VGND sg13g2_decap_8
X_3065_ VGND VPWR _0853_ _0855_ tmds_red.n114 tmds_red.n100 sg13g2_a21oi_2
X_4981__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_23_402 VPWR VGND sg13g2_fill_1
XFILLER_24_925 VPWR VGND sg13g2_decap_8
XFILLER_23_435 VPWR VGND sg13g2_decap_8
X_3967_ _1658_ VPWR _1693_ VGND _1673_ _1691_ sg13g2_o21ai_1
X_2918_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\] net753 _0788_ _0286_
+ VPWR VGND sg13g2_mux2_1
X_3898_ _1623_ VPWR _1624_ VGND _1174_ _1622_ sg13g2_o21ai_1
X_2849_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\] _0774_ _0415_
+ VPWR VGND sg13g2_mux2_1
XFILLER_2_306 VPWR VGND sg13g2_fill_2
X_4519_ net676 net728 _0072_ VPWR VGND sg13g2_nor2_1
XFILLER_5_8 VPWR VGND sg13g2_fill_2
Xfanout610 videogen.fancy_shader.n646\[8\] net610 VPWR VGND sg13g2_buf_8
Xfanout632 net650 net632 VPWR VGND sg13g2_buf_8
Xfanout621 net623 net621 VPWR VGND sg13g2_buf_8
Xfanout665 net667 net665 VPWR VGND sg13g2_buf_1
Xfanout676 net678 net676 VPWR VGND sg13g2_buf_8
Xfanout654 net655 net654 VPWR VGND sg13g2_buf_1
Xfanout643 net650 net643 VPWR VGND sg13g2_buf_8
Xfanout698 net701 net698 VPWR VGND sg13g2_buf_2
Xfanout687 net693 net687 VPWR VGND sg13g2_buf_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_19_719 VPWR VGND sg13g2_decap_8
XFILLER_2_1000 VPWR VGND sg13g2_decap_8
X_4960__379 VPWR VGND net379 sg13g2_tiehi
XFILLER_27_774 VPWR VGND sg13g2_decap_8
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_4
XFILLER_6_612 VPWR VGND sg13g2_decap_8
XFILLER_5_122 VPWR VGND sg13g2_decap_8
XFILLER_5_133 VPWR VGND sg13g2_fill_2
XFILLER_6_689 VPWR VGND sg13g2_fill_1
XFILLER_45_9 VPWR VGND sg13g2_fill_1
XFILLER_5_199 VPWR VGND sg13g2_decap_4
XFILLER_49_310 VPWR VGND sg13g2_decap_8
XFILLER_2_895 VPWR VGND sg13g2_decap_8
XFILLER_49_387 VPWR VGND sg13g2_decap_8
XFILLER_37_538 VPWR VGND sg13g2_decap_8
XFILLER_45_571 VPWR VGND sg13g2_fill_2
X_4870_ net259 VGND VPWR _0421_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\]
+ _0078_ sg13g2_dfrbpq_1
X_3821_ _1551_ _1450_ _1549_ _1251_ _1250_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_276 VPWR VGND sg13g2_fill_1
X_3752_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\] net559 _1482_ VPWR
+ VGND sg13g2_nor2_1
X_3683_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\] net549 _1413_ VPWR
+ VGND sg13g2_nor2_1
X_2703_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\] _0740_ _0536_
+ VPWR VGND sg13g2_mux2_1
X_2634_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\] net774 _0722_ _0587_
+ VPWR VGND sg13g2_mux2_1
X_2565_ _0680_ net543 _0678_ VPWR VGND sg13g2_nand2_2
X_4304_ net606 VPWR _2005_ VGND _2002_ _2004_ sg13g2_o21ai_1
XFILLER_4_70 VPWR VGND sg13g2_decap_4
X_4235_ _1941_ _1932_ _1942_ VPWR VGND sg13g2_xor2_1
X_4166_ net1 VPWR _1889_ VGND _1880_ _1888_ sg13g2_o21ai_1
X_3117_ net751 _0795_ _0900_ _0305_ VPWR VGND sg13g2_nor3_1
XFILLER_28_516 VPWR VGND sg13g2_fill_2
X_4097_ _1819_ _1120_ _1820_ VPWR VGND sg13g2_xor2_1
X_3048_ tmds_green.dc_balancing_reg\[0\] tmds_green.dc_balancing_reg\[1\] tmds_green.dc_balancing_reg\[3\]
+ tmds_green.dc_balancing_reg\[2\] _0839_ VPWR VGND sg13g2_nor4_1
X_4840__317 VPWR VGND net317 sg13g2_tiehi
XFILLER_24_733 VPWR VGND sg13g2_decap_8
XFILLER_12_939 VPWR VGND sg13g2_decap_8
X_4999_ net199 VGND VPWR _0546_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\]
+ _0194_ sg13g2_dfrbpq_1
XFILLER_2_103 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_24_1023 VPWR VGND sg13g2_decap_4
XFILLER_48_87 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_27_593 VPWR VGND sg13g2_decap_8
XFILLER_30_703 VPWR VGND sg13g2_decap_8
XFILLER_30_747 VPWR VGND sg13g2_fill_1
XFILLER_30_769 VPWR VGND sg13g2_decap_4
XFILLER_7_954 VPWR VGND sg13g2_decap_8
XFILLER_6_453 VPWR VGND sg13g2_fill_1
XFILLER_2_681 VPWR VGND sg13g2_decap_4
X_4020_ VGND VPWR _1739_ _1741_ _1743_ _1736_ sg13g2_a21oi_1
XFILLER_1_180 VPWR VGND sg13g2_decap_8
XFILLER_37_302 VPWR VGND sg13g2_decap_8
XFILLER_49_195 VPWR VGND sg13g2_decap_8
XFILLER_38_858 VPWR VGND sg13g2_fill_1
X_4922_ net144 VGND VPWR _0473_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\]
+ _0130_ sg13g2_dfrbpq_1
XFILLER_21_703 VPWR VGND sg13g2_decap_8
X_4853_ net292 VGND VPWR _0404_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\]
+ _0061_ sg13g2_dfrbpq_1
XFILLER_21_725 VPWR VGND sg13g2_decap_8
X_4784_ net34 VGND VPWR _0335_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ net633 sg13g2_dfrbpq_1
XFILLER_20_246 VPWR VGND sg13g2_decap_8
X_3804_ net617 VPWR _1534_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\]
+ net577 sg13g2_o21ai_1
X_3735_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\] net584 _1465_ VPWR
+ VGND sg13g2_nor2_1
X_3666_ _1392_ _1393_ _1394_ _1395_ _1396_ VPWR VGND sg13g2_nor4_1
Xheichips25_bagel_28 VPWR VGND uio_oe[7] sg13g2_tielo
X_3597_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\] net584 _1327_ VPWR
+ VGND sg13g2_nor2_1
X_2617_ _0716_ _0713_ _0715_ VPWR VGND sg13g2_nand2_2
XFILLER_0_618 VPWR VGND sg13g2_decap_8
X_2548_ net608 net609 _0663_ VPWR VGND sg13g2_nor2_1
X_4218_ VGND VPWR _0843_ _1927_ _0500_ net750 sg13g2_a21oi_1
XFILLER_29_803 VPWR VGND sg13g2_decap_8
XFILLER_18_24 VPWR VGND sg13g2_fill_1
XFILLER_28_324 VPWR VGND sg13g2_fill_1
X_4149_ _1870_ _1871_ _1872_ VPWR VGND sg13g2_nor2_1
XFILLER_43_338 VPWR VGND sg13g2_decap_8
XFILLER_43_327 VPWR VGND sg13g2_fill_1
XFILLER_37_891 VPWR VGND sg13g2_decap_4
XFILLER_11_213 VPWR VGND sg13g2_fill_2
XFILLER_24_585 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_fill_2
Xclkload0 VPWR clkload0/Y clknet_1_1__leaf_clk VGND sg13g2_inv_1
XFILLER_4_957 VPWR VGND sg13g2_decap_8
XFILLER_47_611 VPWR VGND sg13g2_decap_8
XFILLER_46_121 VPWR VGND sg13g2_fill_2
XFILLER_35_817 VPWR VGND sg13g2_decap_4
XFILLER_34_349 VPWR VGND sg13g2_decap_4
XFILLER_27_390 VPWR VGND sg13g2_decap_4
XFILLER_30_500 VPWR VGND sg13g2_fill_1
XFILLER_30_533 VPWR VGND sg13g2_decap_8
XFILLER_30_544 VPWR VGND sg13g2_fill_2
X_3520_ _1249_ _1248_ _1241_ _1250_ VPWR VGND sg13g2_a21o_2
XFILLER_7_795 VPWR VGND sg13g2_fill_2
X_3451_ _1158_ net547 _1181_ VPWR VGND sg13g2_nor2_1
X_3382_ _1112_ _1099_ _1110_ VPWR VGND sg13g2_xnor2_1
X_5121_ net799 VGND VPWR serialize.n427\[5\] serialize.n411\[3\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5052_ net72 VGND VPWR _0599_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\]
+ _0247_ sg13g2_dfrbpq_1
XFILLER_38_622 VPWR VGND sg13g2_decap_4
X_4003_ _1039_ _1725_ _1726_ VPWR VGND sg13g2_nor2_2
XFILLER_26_806 VPWR VGND sg13g2_fill_1
XFILLER_1_82 VPWR VGND sg13g2_decap_4
XFILLER_34_872 VPWR VGND sg13g2_fill_2
X_4904__188 VPWR VGND net188 sg13g2_tiehi
X_4905_ net186 VGND VPWR _0456_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\]
+ _0113_ sg13g2_dfrbpq_1
X_4836_ net323 VGND VPWR _0387_ red_tmds_par\[8\] net642 sg13g2_dfrbpq_1
XFILLER_21_588 VPWR VGND sg13g2_decap_4
X_4767_ net68 VGND VPWR _0318_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\]
+ net631 sg13g2_dfrbpq_2
X_4698_ net690 net744 _0251_ VPWR VGND sg13g2_nor2_1
XFILLER_4_209 VPWR VGND sg13g2_decap_8
X_3718_ _0650_ _1447_ _1448_ VPWR VGND sg13g2_nor2_1
X_3649_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\] net572 _1379_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_36 VPWR VGND sg13g2_fill_2
XFILLER_1_916 VPWR VGND sg13g2_decap_8
Xhold12 serialize.n414\[1\] VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold23 serialize.n428\[6\] VPWR VGND net428 sg13g2_dlygate4sd3_1
XFILLER_0_448 VPWR VGND sg13g2_fill_2
Xhold34 serialize.n414\[7\] VPWR VGND net439 sg13g2_dlygate4sd3_1
XFILLER_29_78 VPWR VGND sg13g2_decap_8
XFILLER_29_600 VPWR VGND sg13g2_decap_4
XFILLER_29_611 VPWR VGND sg13g2_fill_1
XFILLER_45_22 VPWR VGND sg13g2_decap_4
XFILLER_31_319 VPWR VGND sg13g2_fill_2
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_24_393 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_fill_2
XFILLER_12_577 VPWR VGND sg13g2_decap_8
XFILLER_6_27 VPWR VGND sg13g2_decap_8
XFILLER_0_982 VPWR VGND sg13g2_decap_8
XFILLER_19_110 VPWR VGND sg13g2_fill_1
XFILLER_48_986 VPWR VGND sg13g2_decap_8
XFILLER_19_143 VPWR VGND sg13g2_decap_4
XFILLER_34_102 VPWR VGND sg13g2_fill_1
XFILLER_16_850 VPWR VGND sg13g2_fill_1
XFILLER_35_658 VPWR VGND sg13g2_fill_1
XFILLER_37_1011 VPWR VGND sg13g2_decap_8
X_2951_ VGND VPWR _0809_ videogen.test_lut_thingy.pixel_feeder_inst.state\[3\] videogen.test_lut_thingy.pixel_feeder_inst.state\[1\]
+ sg13g2_or2_1
XFILLER_43_691 VPWR VGND sg13g2_decap_4
X_2882_ _0689_ _0725_ _0781_ VPWR VGND sg13g2_nor2_2
X_4621_ net688 net742 _0174_ VPWR VGND sg13g2_nor2_1
X_4552_ net680 net731 _0105_ VPWR VGND sg13g2_nor2_1
X_4483_ net670 net721 _0036_ VPWR VGND sg13g2_nor2_1
X_3503_ _1226_ VPWR _1233_ VGND _1227_ _1232_ sg13g2_o21ai_1
X_3434_ _1164_ _1162_ _1163_ VPWR VGND sg13g2_nand2_1
X_3365_ videogen.fancy_shader.video_y\[8\] net610 _1095_ VPWR VGND sg13g2_nor2_1
X_5104_ net800 VGND VPWR serialize.n429\[1\] serialize.n458 clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3296_ _1015_ _1017_ _1026_ VPWR VGND sg13g2_and2_1
X_5035_ net264 VGND VPWR _0582_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\]
+ _0230_ sg13g2_dfrbpq_1
XFILLER_39_986 VPWR VGND sg13g2_decap_8
XFILLER_26_636 VPWR VGND sg13g2_decap_8
XFILLER_25_135 VPWR VGND sg13g2_decap_8
XFILLER_25_146 VPWR VGND sg13g2_decap_4
XFILLER_41_639 VPWR VGND sg13g2_decap_4
XFILLER_41_617 VPWR VGND sg13g2_fill_1
X_4806__362 VPWR VGND net362 sg13g2_tiehi
XFILLER_25_168 VPWR VGND sg13g2_decap_4
XFILLER_40_149 VPWR VGND sg13g2_decap_4
XFILLER_22_831 VPWR VGND sg13g2_decap_8
XFILLER_21_352 VPWR VGND sg13g2_decap_4
XFILLER_22_886 VPWR VGND sg13g2_decap_8
X_4991__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_21_396 VPWR VGND sg13g2_decap_8
X_4819_ net340 VGND VPWR _0370_ hsync net640 sg13g2_dfrbpq_2
XFILLER_5_529 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_212 VPWR VGND sg13g2_decap_8
XFILLER_1_713 VPWR VGND sg13g2_decap_8
XFILLER_0_256 VPWR VGND sg13g2_decap_8
XFILLER_45_901 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk_regs clknet_0_clk_regs clknet_3_0__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_29_463 VPWR VGND sg13g2_fill_1
XFILLER_45_978 VPWR VGND sg13g2_decap_8
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_32_639 VPWR VGND sg13g2_decap_8
XFILLER_12_363 VPWR VGND sg13g2_fill_1
X_3150_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0922_ _0923_ VPWR VGND
+ sg13g2_and2_1
XFILLER_39_249 VPWR VGND sg13g2_fill_1
XFILLER_39_238 VPWR VGND sg13g2_fill_2
X_3081_ _0871_ _0859_ _0869_ VPWR VGND sg13g2_xnor2_1
X_4788__398 VPWR VGND net398 sg13g2_tiehi
XFILLER_22_116 VPWR VGND sg13g2_decap_8
X_3983_ _1701_ _1704_ _1625_ _1709_ VPWR VGND sg13g2_nand3_1
X_2934_ net793 _0792_ _0371_ VPWR VGND sg13g2_and2_1
XFILLER_31_661 VPWR VGND sg13g2_decap_8
X_2865_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\] net773 _0777_ _0402_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_160 VPWR VGND sg13g2_decap_8
X_4604_ net666 net717 _0157_ VPWR VGND sg13g2_nor2_1
X_4535_ net659 net710 _0088_ VPWR VGND sg13g2_nor2_1
X_2796_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\] _0759_ _0453_
+ VPWR VGND sg13g2_mux2_1
X_4871__257 VPWR VGND net257 sg13g2_tiehi
X_4466_ net674 net725 _0019_ VPWR VGND sg13g2_nor2_1
X_4397_ _2088_ _2074_ _2086_ VPWR VGND sg13g2_xnor2_1
X_3417_ VGND VPWR _1147_ _1146_ _1145_ sg13g2_or2_1
Xfanout803 rst_n net803 VPWR VGND sg13g2_buf_8
X_3348_ _1050_ VPWR _1078_ VGND _0633_ _0634_ sg13g2_o21ai_1
X_3279_ videogen.fancy_shader.n646\[2\] videogen.fancy_shader.video_y\[2\] _1009_
+ VPWR VGND sg13g2_xor2_1
XFILLER_27_912 VPWR VGND sg13g2_decap_8
XFILLER_38_260 VPWR VGND sg13g2_decap_4
X_5018_ net67 VGND VPWR _0565_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\]
+ _0213_ sg13g2_dfrbpq_1
XFILLER_26_433 VPWR VGND sg13g2_fill_2
XFILLER_27_989 VPWR VGND sg13g2_decap_8
XFILLER_42_937 VPWR VGND sg13g2_decap_8
XFILLER_26_68 VPWR VGND sg13g2_decap_8
XFILLER_13_149 VPWR VGND sg13g2_decap_8
XFILLER_42_34 VPWR VGND sg13g2_decap_8
XFILLER_41_469 VPWR VGND sg13g2_decap_4
XFILLER_10_856 VPWR VGND sg13g2_fill_1
XFILLER_5_359 VPWR VGND sg13g2_decap_8
XFILLER_27_1010 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_18_945 VPWR VGND sg13g2_decap_8
XFILLER_36_219 VPWR VGND sg13g2_decap_8
XFILLER_17_433 VPWR VGND sg13g2_decap_4
XFILLER_17_477 VPWR VGND sg13g2_decap_8
XFILLER_32_469 VPWR VGND sg13g2_decap_4
XFILLER_34_1014 VPWR VGND sg13g2_decap_8
X_2650_ _0729_ _0713_ _0727_ VPWR VGND sg13g2_nand2_2
XFILLER_8_131 VPWR VGND sg13g2_decap_8
X_2581_ _0692_ _0695_ _0696_ VPWR VGND sg13g2_nor2_1
X_4320_ _2015_ _2016_ net602 _2017_ VPWR VGND sg13g2_nand3_1
X_4251_ _1956_ _1955_ _1957_ VPWR VGND sg13g2_xor2_1
X_3202_ _0635_ _0918_ _0957_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1007 VPWR VGND sg13g2_decap_8
X_4182_ _1352_ _1720_ _1904_ VPWR VGND sg13g2_nor2_1
X_3133_ _0908_ videogen.fancy_shader.video_x\[9\] _0910_ VPWR VGND sg13g2_xor2_1
XFILLER_28_709 VPWR VGND sg13g2_decap_8
XFILLER_27_219 VPWR VGND sg13g2_decap_8
X_3064_ _0854_ tmds_red.n126 tmds_red.n132 VPWR VGND sg13g2_xnor2_1
XFILLER_24_904 VPWR VGND sg13g2_decap_8
X_3966_ _1657_ _1672_ _1692_ VPWR VGND _1691_ sg13g2_nand3b_1
X_2917_ _0699_ _0721_ _0788_ VPWR VGND sg13g2_nor2_2
X_3897_ _1623_ _1006_ _1622_ VPWR VGND sg13g2_nand2_2
X_2848_ net756 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\] _0774_ _0416_
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_37 VPWR VGND sg13g2_decap_4
X_2779_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\] _0756_ _0467_
+ VPWR VGND sg13g2_mux2_1
X_4518_ net674 net726 _0071_ VPWR VGND sg13g2_nor2_1
XFILLER_2_329 VPWR VGND sg13g2_fill_1
X_4449_ _1989_ VPWR _2138_ VGND _2135_ _2137_ sg13g2_o21ai_1
Xfanout633 net634 net633 VPWR VGND sg13g2_buf_8
Xfanout600 videogen.mem_read net600 VPWR VGND sg13g2_buf_8
Xfanout611 videogen.fancy_shader.n646\[3\] net611 VPWR VGND sg13g2_buf_8
Xfanout622 net623 net622 VPWR VGND sg13g2_buf_8
Xfanout666 net667 net666 VPWR VGND sg13g2_buf_8
Xfanout644 net646 net644 VPWR VGND sg13g2_buf_8
Xfanout655 net656 net655 VPWR VGND sg13g2_buf_8
Xfanout699 net701 net699 VPWR VGND sg13g2_buf_8
Xfanout677 net678 net677 VPWR VGND sg13g2_buf_1
Xfanout688 net689 net688 VPWR VGND sg13g2_buf_8
XFILLER_46_517 VPWR VGND sg13g2_fill_1
XFILLER_37_67 VPWR VGND sg13g2_fill_2
XFILLER_27_786 VPWR VGND sg13g2_fill_2
XFILLER_41_222 VPWR VGND sg13g2_decap_8
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_42_789 VPWR VGND sg13g2_decap_4
XFILLER_41_288 VPWR VGND sg13g2_fill_1
XFILLER_10_631 VPWR VGND sg13g2_fill_1
XFILLER_10_653 VPWR VGND sg13g2_decap_8
XFILLER_5_101 VPWR VGND sg13g2_decap_8
XFILLER_10_686 VPWR VGND sg13g2_fill_2
XFILLER_2_874 VPWR VGND sg13g2_decap_8
XFILLER_49_366 VPWR VGND sg13g2_decap_8
XFILLER_33_734 VPWR VGND sg13g2_fill_2
XFILLER_21_929 VPWR VGND sg13g2_decap_8
X_3820_ VPWR _1550_ _1549_ VGND sg13g2_inv_1
XFILLER_32_244 VPWR VGND sg13g2_fill_1
X_3751_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\] net572 _1481_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_14_992 VPWR VGND sg13g2_decap_8
X_2702_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\] _0740_ _0537_
+ VPWR VGND sg13g2_mux2_1
X_3682_ net614 VPWR _1412_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[1\]
+ net572 sg13g2_o21ai_1
X_4781__40 VPWR VGND net40 sg13g2_tiehi
X_2633_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\] net764 _0722_ _0588_
+ VPWR VGND sg13g2_mux2_1
X_2564_ net543 _0678_ _0679_ VPWR VGND sg13g2_and2_1
X_4303_ net604 _1989_ _2004_ VPWR VGND sg13g2_nor2_2
X_4234_ _1934_ _1935_ _1941_ VPWR VGND sg13g2_nor2_1
X_4165_ _1887_ _1879_ _1888_ VPWR VGND sg13g2_nor2b_1
X_3116_ VGND VPWR videogen.fancy_shader.video_x\[1\] net630 _0900_ videogen.fancy_shader.video_x\[2\]
+ sg13g2_a21oi_1
X_4096_ _1819_ _1730_ _1807_ VPWR VGND sg13g2_xnor2_1
X_3047_ _0642_ net569 _0271_ VPWR VGND sg13g2_nor2_1
XFILLER_24_712 VPWR VGND sg13g2_decap_8
XFILLER_36_594 VPWR VGND sg13g2_fill_2
XFILLER_12_918 VPWR VGND sg13g2_decap_8
XFILLER_24_756 VPWR VGND sg13g2_fill_1
X_4998_ net203 VGND VPWR _0545_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\]
+ _0193_ sg13g2_dfrbpq_1
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_23_299 VPWR VGND sg13g2_fill_1
X_4877__241 VPWR VGND net241 sg13g2_tiehi
X_3949_ _1675_ _1672_ _1674_ VPWR VGND sg13g2_nand2_1
XFILLER_23_69 VPWR VGND sg13g2_decap_8
XFILLER_20_984 VPWR VGND sg13g2_decap_8
XFILLER_2_115 VPWR VGND sg13g2_decap_8
X_4914__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
XFILLER_19_539 VPWR VGND sg13g2_fill_1
XFILLER_46_369 VPWR VGND sg13g2_decap_8
XFILLER_27_572 VPWR VGND sg13g2_decap_8
XFILLER_14_200 VPWR VGND sg13g2_fill_2
XFILLER_14_233 VPWR VGND sg13g2_decap_8
XFILLER_14_255 VPWR VGND sg13g2_decap_8
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_6_465 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_fill_1
XFILLER_49_141 VPWR VGND sg13g2_decap_8
XFILLER_29_5 VPWR VGND sg13g2_fill_2
XFILLER_49_174 VPWR VGND sg13g2_decap_8
X_4921_ net148 VGND VPWR _0472_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\]
+ _0129_ sg13g2_dfrbpq_1
X_4852_ net294 VGND VPWR _0403_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\]
+ _0060_ sg13g2_dfrbpq_1
X_3803_ net594 _1527_ _1532_ _1533_ VPWR VGND sg13g2_nor3_1
X_4783_ net36 VGND VPWR _0334_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\]
+ net633 sg13g2_dfrbpq_1
X_3734_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\] net551 _1464_ VPWR
+ VGND sg13g2_nor2_1
X_3665_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\] net584 _1395_ VPWR
+ VGND sg13g2_nor2_1
Xheichips25_bagel_29 VPWR VGND uio_out[1] sg13g2_tielo
X_2616_ _0715_ net592 _0692_ _0697_ VPWR VGND sg13g2_and3_2
X_3596_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\] net574 _1326_ VPWR
+ VGND sg13g2_nor2_1
X_2547_ _0662_ _0661_ videogen.fancy_shader.video_y\[4\] VPWR VGND sg13g2_nand2b_1
X_4217_ net607 _0846_ _1927_ VPWR VGND sg13g2_and2_1
X_4148_ _1871_ _1798_ _1866_ _1869_ VPWR VGND sg13g2_and3_1
XFILLER_29_848 VPWR VGND sg13g2_fill_2
XFILLER_43_306 VPWR VGND sg13g2_fill_2
X_4079_ _1802_ _1055_ _1800_ VPWR VGND sg13g2_xnor2_1
X_5044__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_24_553 VPWR VGND sg13g2_decap_8
XFILLER_8_708 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_3_0__leaf_clk_regs clkload1/X VPWR VGND sg13g2_buf_1
XFILLER_4_936 VPWR VGND sg13g2_decap_8
XFILLER_3_446 VPWR VGND sg13g2_decap_8
XFILLER_34_306 VPWR VGND sg13g2_fill_2
XFILLER_15_553 VPWR VGND sg13g2_fill_2
XFILLER_15_597 VPWR VGND sg13g2_fill_2
XFILLER_30_578 VPWR VGND sg13g2_decap_8
XFILLER_7_752 VPWR VGND sg13g2_decap_8
XFILLER_11_792 VPWR VGND sg13g2_decap_8
XFILLER_6_262 VPWR VGND sg13g2_decap_4
XFILLER_6_295 VPWR VGND sg13g2_fill_1
X_3450_ _1173_ net547 _1180_ VPWR VGND sg13g2_nor2_1
X_3381_ _1110_ _1099_ _1111_ VPWR VGND sg13g2_xor2_1
X_5120_ net798 VGND VPWR serialize.n427\[4\] serialize.n411\[2\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5051_ net98 VGND VPWR _0598_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\]
+ _0246_ sg13g2_dfrbpq_1
X_4002_ VGND VPWR _1725_ _1724_ _1013_ sg13g2_or2_1
XFILLER_38_678 VPWR VGND sg13g2_decap_4
XFILLER_25_328 VPWR VGND sg13g2_decap_8
XFILLER_34_851 VPWR VGND sg13g2_decap_8
X_4904_ net188 VGND VPWR _0455_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\]
+ _0112_ sg13g2_dfrbpq_1
X_4835_ net324 VGND VPWR _0386_ red_tmds_par\[6\] net644 sg13g2_dfrbpq_1
XFILLER_21_567 VPWR VGND sg13g2_decap_8
X_4798__378 VPWR VGND net378 sg13g2_tiehi
X_4766_ net69 VGND VPWR _0317_ tmds_blue.vsync net640 sg13g2_dfrbpq_1
X_3717_ _0636_ _1423_ _1446_ _1447_ VPWR VGND sg13g2_nor3_1
X_4697_ net690 net744 _0250_ VPWR VGND sg13g2_nor2_1
X_3648_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\] net559 _1378_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_48 VPWR VGND sg13g2_decap_8
X_3579_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\] net588 _1309_ VPWR
+ VGND sg13g2_nor2_1
Xhold13 serialize.n417\[6\] VPWR VGND net418 sg13g2_dlygate4sd3_1
XFILLER_48_409 VPWR VGND sg13g2_fill_1
Xhold24 serialize.bit_cnt\[1\] VPWR VGND net429 sg13g2_dlygate4sd3_1
Xhold35 serialize.n414\[2\] VPWR VGND net440 sg13g2_dlygate4sd3_1
XFILLER_29_57 VPWR VGND sg13g2_decap_8
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_100 VPWR VGND sg13g2_decap_8
XFILLER_29_645 VPWR VGND sg13g2_fill_2
XFILLER_29_656 VPWR VGND sg13g2_fill_2
X_4729__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_45_45 VPWR VGND sg13g2_decap_8
XFILLER_45_34 VPWR VGND sg13g2_fill_1
XFILLER_45_67 VPWR VGND sg13g2_fill_2
XFILLER_6_39 VPWR VGND sg13g2_decap_4
XFILLER_4_744 VPWR VGND sg13g2_fill_2
XFILLER_4_722 VPWR VGND sg13g2_decap_8
XFILLER_0_961 VPWR VGND sg13g2_decap_8
XFILLER_13_8 VPWR VGND sg13g2_decap_4
XFILLER_48_965 VPWR VGND sg13g2_decap_8
XFILLER_34_114 VPWR VGND sg13g2_fill_1
XFILLER_35_637 VPWR VGND sg13g2_fill_1
X_2950_ _0808_ videogen.test_lut_thingy.pixel_feeder_inst.state\[1\] _0792_ VPWR VGND
+ sg13g2_nand2b_1
XFILLER_15_361 VPWR VGND sg13g2_decap_8
X_2881_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\] net783 _0780_ _0389_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_383 VPWR VGND sg13g2_decap_8
XFILLER_31_832 VPWR VGND sg13g2_fill_1
X_4620_ net692 net741 _0173_ VPWR VGND sg13g2_nor2_1
X_4551_ net680 net730 _0104_ VPWR VGND sg13g2_nor2_1
X_4482_ net670 net721 _0035_ VPWR VGND sg13g2_nor2_1
X_3502_ net547 VPWR _1232_ VGND _1228_ _1231_ sg13g2_o21ai_1
X_3433_ _1134_ _1145_ _1161_ _1163_ VPWR VGND sg13g2_or3_1
X_5103_ net800 VGND VPWR serialize.n429\[0\] serialize.n456 clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_3364_ VPWR VGND _1080_ _1090_ _1093_ _1081_ _1094_ _1091_ sg13g2_a221oi_1
XFILLER_32_0 VPWR VGND sg13g2_fill_1
X_3295_ videogen.fancy_shader.video_x\[3\] net611 _1025_ VPWR VGND sg13g2_xor2_1
X_5034_ net271 VGND VPWR _0581_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\]
+ _0229_ sg13g2_dfrbpq_1
XFILLER_39_965 VPWR VGND sg13g2_decap_8
XFILLER_38_464 VPWR VGND sg13g2_fill_2
XFILLER_15_26 VPWR VGND sg13g2_fill_1
XFILLER_22_810 VPWR VGND sg13g2_decap_8
XFILLER_22_865 VPWR VGND sg13g2_decap_8
XFILLER_33_191 VPWR VGND sg13g2_fill_1
X_4818_ net341 VGND VPWR _0369_ videogen.test_lut_thingy.gol_counter_reg\[3\] net643
+ sg13g2_dfrbpq_1
X_4749_ net93 VGND VPWR _0300_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\]
+ _0031_ sg13g2_dfrbpq_1
Xoutput14 net14 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_769 VPWR VGND sg13g2_decap_8
XFILLER_48_206 VPWR VGND sg13g2_decap_4
XFILLER_48_239 VPWR VGND sg13g2_decap_4
X_4963__367 VPWR VGND net367 sg13g2_tiehi
XFILLER_44_412 VPWR VGND sg13g2_fill_2
XFILLER_45_957 VPWR VGND sg13g2_decap_8
XFILLER_16_136 VPWR VGND sg13g2_fill_1
XFILLER_40_651 VPWR VGND sg13g2_decap_8
X_4970__316 VPWR VGND net316 sg13g2_tiehi
X_3080_ _0870_ _0861_ _0869_ VPWR VGND sg13g2_nand2_1
XFILLER_48_740 VPWR VGND sg13g2_decap_8
X_4829__330 VPWR VGND net330 sg13g2_tiehi
XFILLER_36_946 VPWR VGND sg13g2_decap_8
XFILLER_35_445 VPWR VGND sg13g2_decap_8
XFILLER_36_957 VPWR VGND sg13g2_fill_2
X_3982_ _1698_ _1707_ _1708_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_618 VPWR VGND sg13g2_decap_8
X_2933_ videogen.fancy_shader.video_y\[9\] _0661_ _0667_ _0792_ VGND VPWR _0791_ sg13g2_nor4_2
X_5052__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_15_191 VPWR VGND sg13g2_fill_1
XFILLER_31_640 VPWR VGND sg13g2_decap_4
X_2864_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\] net764 _0777_ _0403_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_695 VPWR VGND sg13g2_fill_1
X_2795_ net778 videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\] _0759_ _0454_
+ VPWR VGND sg13g2_mux2_1
X_4603_ net668 net720 _0156_ VPWR VGND sg13g2_nor2_1
XFILLER_8_891 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
X_4534_ net660 net711 _0087_ VPWR VGND sg13g2_nor2_1
X_4836__323 VPWR VGND net323 sg13g2_tiehi
X_4465_ net675 net725 _0018_ VPWR VGND sg13g2_nor2_1
X_4396_ _2074_ _2086_ _2087_ VPWR VGND sg13g2_and2_1
X_3416_ net544 _1140_ _1144_ _1146_ VPWR VGND sg13g2_nor3_1
X_3347_ VGND VPWR _1077_ _1061_ _1051_ sg13g2_or2_1
XFILLER_45_209 VPWR VGND sg13g2_decap_4
XFILLER_39_762 VPWR VGND sg13g2_decap_8
X_3278_ videogen.fancy_shader.video_y\[2\] videogen.fancy_shader.n646\[2\] _1008_
+ VPWR VGND sg13g2_and2_1
X_5017_ net76 VGND VPWR _0564_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\]
+ _0212_ sg13g2_dfrbpq_1
XFILLER_27_968 VPWR VGND sg13g2_decap_8
XFILLER_42_916 VPWR VGND sg13g2_decap_8
XFILLER_14_618 VPWR VGND sg13g2_decap_4
XFILLER_26_478 VPWR VGND sg13g2_decap_8
XFILLER_42_79 VPWR VGND sg13g2_fill_2
XFILLER_10_879 VPWR VGND sg13g2_fill_2
XFILLER_49_504 VPWR VGND sg13g2_decap_8
XFILLER_18_924 VPWR VGND sg13g2_decap_8
XFILLER_29_250 VPWR VGND sg13g2_fill_1
XFILLER_44_253 VPWR VGND sg13g2_fill_2
XFILLER_41_993 VPWR VGND sg13g2_decap_8
XFILLER_9_633 VPWR VGND sg13g2_fill_1
XFILLER_12_172 VPWR VGND sg13g2_decap_4
XFILLER_13_673 VPWR VGND sg13g2_decap_8
XFILLER_8_198 VPWR VGND sg13g2_decap_8
X_2580_ net543 _0694_ _0695_ VPWR VGND sg13g2_and2_1
XFILLER_5_883 VPWR VGND sg13g2_decap_8
XFILLER_4_393 VPWR VGND sg13g2_decap_8
X_4250_ VGND VPWR _0654_ _0883_ _1956_ _0886_ sg13g2_a21oi_1
X_3201_ _0951_ _0956_ _0337_ VPWR VGND sg13g2_nor2_1
X_4181_ VGND VPWR _1900_ _1903_ _0381_ net750 sg13g2_a21oi_1
X_3132_ _0898_ _0909_ _0311_ VPWR VGND sg13g2_nor2_1
X_3063_ _0850_ _0851_ _0852_ _0853_ VPWR VGND sg13g2_nor3_1
XFILLER_35_231 VPWR VGND sg13g2_fill_2
X_3965_ VPWR VGND _1683_ _1675_ _1671_ _1627_ _1691_ _1628_ sg13g2_a221oi_1
XFILLER_23_459 VPWR VGND sg13g2_fill_1
X_2916_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\] net787 _0787_ _0287_
+ VPWR VGND sg13g2_mux2_1
X_3896_ videogen.fancy_shader.n646\[0\] videogen.fancy_shader.video_y\[0\] _1622_
+ VPWR VGND sg13g2_xor2_1
XFILLER_12_16 VPWR VGND sg13g2_decap_8
X_2847_ _0774_ _0710_ _0773_ VPWR VGND sg13g2_nand2_2
XFILLER_31_481 VPWR VGND sg13g2_fill_2
X_2778_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\] _0756_ _0468_
+ VPWR VGND sg13g2_mux2_1
X_4517_ net675 net725 _0070_ VPWR VGND sg13g2_nor2_1
XFILLER_2_308 VPWR VGND sg13g2_fill_1
X_4448_ _2123_ _2136_ _2137_ VPWR VGND _1991_ sg13g2_nand3b_1
Xfanout623 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\] net623 VPWR VGND
+ sg13g2_buf_8
Xfanout612 net613 net612 VPWR VGND sg13g2_buf_8
Xfanout601 tmds_green.n132 net601 VPWR VGND sg13g2_buf_8
Xfanout667 net673 net667 VPWR VGND sg13g2_buf_8
X_4379_ VGND VPWR _2063_ _2072_ _0622_ net570 sg13g2_a21oi_1
Xfanout645 net646 net645 VPWR VGND sg13g2_buf_1
Xfanout634 net635 net634 VPWR VGND sg13g2_buf_8
Xfanout656 net694 net656 VPWR VGND sg13g2_buf_8
XFILLER_46_507 VPWR VGND sg13g2_decap_4
X_5047__165 VPWR VGND net165 sg13g2_tiehi
Xfanout678 net683 net678 VPWR VGND sg13g2_buf_8
Xfanout689 net692 net689 VPWR VGND sg13g2_buf_8
XFILLER_46_529 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_4
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_fill_1
XFILLER_41_267 VPWR VGND sg13g2_decap_8
X_5016__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_6_647 VPWR VGND sg13g2_fill_2
XFILLER_5_146 VPWR VGND sg13g2_decap_4
X_4819__340 VPWR VGND net340 sg13g2_tiehi
XFILLER_2_853 VPWR VGND sg13g2_decap_8
XFILLER_49_345 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_fill_2
X_4826__333 VPWR VGND net333 sg13g2_tiehi
XFILLER_45_573 VPWR VGND sg13g2_fill_1
XFILLER_21_908 VPWR VGND sg13g2_decap_8
X_3750_ net614 VPWR _1480_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\]
+ net549 sg13g2_o21ai_1
XFILLER_14_971 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_decap_4
X_2701_ _0740_ _0706_ _0710_ VPWR VGND sg13g2_nand2_2
X_3681_ net621 _1405_ _1410_ _1411_ VPWR VGND sg13g2_nor3_1
X_2632_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\] net754 _0722_ _0589_
+ VPWR VGND sg13g2_mux2_1
X_2563_ _0676_ _0677_ _0678_ VPWR VGND sg13g2_nor2_2
X_4833__326 VPWR VGND net326 sg13g2_tiehi
X_4302_ VPWR _2003_ _2002_ VGND sg13g2_inv_1
X_4233_ _1929_ _1938_ net548 _1940_ VPWR VGND sg13g2_nand3_1
X_4164_ _1876_ _1882_ _1887_ VPWR VGND sg13g2_nor2_1
X_4095_ _1818_ _1111_ _1815_ VPWR VGND sg13g2_xnor2_1
X_3115_ _0898_ _0899_ _0304_ VPWR VGND sg13g2_nor2_1
XFILLER_28_518 VPWR VGND sg13g2_fill_1
XFILLER_49_890 VPWR VGND sg13g2_decap_8
X_3046_ _0266_ net794 net742 net434 VPWR VGND sg13g2_and3_1
XFILLER_36_551 VPWR VGND sg13g2_decap_4
XFILLER_36_584 VPWR VGND sg13g2_fill_1
X_4997_ net207 VGND VPWR _0544_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\]
+ _0192_ sg13g2_dfrbpq_1
X_3948_ _1660_ _1666_ _1669_ _1674_ VPWR VGND sg13g2_or3_1
X_3879_ _1565_ VPWR _1608_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\]
+ net552 sg13g2_o21ai_1
X_4757__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_20_963 VPWR VGND sg13g2_decap_8
XFILLER_3_628 VPWR VGND sg13g2_fill_2
XFILLER_48_56 VPWR VGND sg13g2_fill_1
XFILLER_7_912 VPWR VGND sg13g2_decap_8
X_4739__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_31_1018 VPWR VGND sg13g2_decap_8
XFILLER_6_422 VPWR VGND sg13g2_decap_4
XFILLER_7_989 VPWR VGND sg13g2_decap_8
XFILLER_2_650 VPWR VGND sg13g2_fill_2
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_160 VPWR VGND sg13g2_fill_2
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_38_805 VPWR VGND sg13g2_decap_8
XFILLER_18_551 VPWR VGND sg13g2_decap_8
XFILLER_46_893 VPWR VGND sg13g2_decap_8
X_4920_ net155 VGND VPWR _0471_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\]
+ _0128_ sg13g2_dfrbpq_1
XFILLER_33_510 VPWR VGND sg13g2_decap_4
X_4851_ net296 VGND VPWR _0402_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\]
+ _0059_ sg13g2_dfrbpq_1
X_3802_ _1528_ _1529_ _1530_ _1531_ _1532_ VPWR VGND sg13g2_nor4_1
X_4782_ net38 VGND VPWR _0333_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\]
+ net632 sg13g2_dfrbpq_1
X_3733_ net596 VPWR _1463_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\]
+ net562 sg13g2_o21ai_1
X_3664_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\] net552 _1394_ VPWR
+ VGND sg13g2_nor2_1
X_2615_ VPWR _0714_ _0713_ VGND sg13g2_inv_1
X_4754__85 VPWR VGND net85 sg13g2_tiehi
X_3595_ net593 VPWR _1325_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\]
+ net561 sg13g2_o21ai_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_2546_ _0633_ _0660_ _0661_ VPWR VGND sg13g2_nor2_1
X_4216_ VGND VPWR tmds_green.n100 net606 _0499_ net750 sg13g2_a21oi_1
X_4147_ VGND VPWR _1866_ _1869_ _1870_ _1798_ sg13g2_a21oi_1
XFILLER_18_15 VPWR VGND sg13g2_decap_8
XFILLER_18_59 VPWR VGND sg13g2_fill_2
X_4078_ _1801_ _1052_ _1799_ VPWR VGND sg13g2_nand2_1
X_3029_ net435 red_tmds_par\[4\] net697 serialize.n427\[4\] VPWR VGND sg13g2_mux2_1
Xclkload2 VPWR clkload2/Y clknet_3_1__leaf_clk_regs VGND sg13g2_inv_1
X_4959__383 VPWR VGND net383 sg13g2_tiehi
XFILLER_20_793 VPWR VGND sg13g2_fill_1
XFILLER_4_915 VPWR VGND sg13g2_decap_8
X_4816__343 VPWR VGND net343 sg13g2_tiehi
XFILLER_1_4 VPWR VGND sg13g2_fill_2
XFILLER_19_304 VPWR VGND sg13g2_fill_2
XFILLER_27_370 VPWR VGND sg13g2_decap_8
XFILLER_28_893 VPWR VGND sg13g2_decap_8
X_4823__336 VPWR VGND net336 sg13g2_tiehi
XFILLER_15_587 VPWR VGND sg13g2_decap_4
XFILLER_10_281 VPWR VGND sg13g2_fill_1
XFILLER_7_797 VPWR VGND sg13g2_fill_1
X_3380_ _1110_ _1108_ _1109_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_981 VPWR VGND sg13g2_decap_8
X_4830__329 VPWR VGND net329 sg13g2_tiehi
XFILLER_34_4 VPWR VGND sg13g2_fill_1
X_5050_ net114 VGND VPWR _0597_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\]
+ _0245_ sg13g2_dfrbpq_1
X_4001_ _1724_ videogen.fancy_shader.n646\[0\] videogen.fancy_shader.video_x\[0\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_37_145 VPWR VGND sg13g2_fill_2
X_4903_ net190 VGND VPWR _0454_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\]
+ _0111_ sg13g2_dfrbpq_1
X_5074__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_21_546 VPWR VGND sg13g2_decap_8
X_4834_ net325 VGND VPWR _0385_ red_tmds_par\[4\] net645 sg13g2_dfrbpq_1
X_4765_ net71 VGND VPWR _0316_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\]
+ _0037_ sg13g2_dfrbpq_1
XFILLER_14_1013 VPWR VGND sg13g2_decap_8
X_3716_ net613 _1434_ _1445_ _1446_ VPWR VGND sg13g2_nor3_1
X_4696_ net664 net715 _0249_ VPWR VGND sg13g2_nor2_1
X_3647_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\] net549 _1377_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_38 VPWR VGND sg13g2_fill_1
X_3578_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\] net555 _1308_ VPWR
+ VGND sg13g2_nor2_1
X_5011__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_0_417 VPWR VGND sg13g2_decap_8
X_2529_ net606 _0647_ VPWR VGND sg13g2_inv_4
Xhold14 serialize.n411\[6\] VPWR VGND net419 sg13g2_dlygate4sd3_1
Xhold25 serialize.n410 VPWR VGND net430 sg13g2_dlygate4sd3_1
Xhold36 serialize.n417\[2\] VPWR VGND net441 sg13g2_dlygate4sd3_1
XFILLER_21_1006 VPWR VGND sg13g2_decap_8
XFILLER_29_624 VPWR VGND sg13g2_fill_2
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_25_830 VPWR VGND sg13g2_fill_1
XFILLER_25_885 VPWR VGND sg13g2_decap_8
XFILLER_40_888 VPWR VGND sg13g2_fill_1
XFILLER_8_517 VPWR VGND sg13g2_fill_1
XFILLER_4_701 VPWR VGND sg13g2_fill_1
XFILLER_3_222 VPWR VGND sg13g2_fill_1
XFILLER_3_277 VPWR VGND sg13g2_fill_2
XFILLER_0_940 VPWR VGND sg13g2_decap_8
XFILLER_48_944 VPWR VGND sg13g2_decap_8
XFILLER_47_432 VPWR VGND sg13g2_decap_4
XFILLER_16_830 VPWR VGND sg13g2_fill_1
XFILLER_35_649 VPWR VGND sg13g2_decap_8
XFILLER_15_340 VPWR VGND sg13g2_decap_8
XFILLER_16_874 VPWR VGND sg13g2_decap_8
XFILLER_31_811 VPWR VGND sg13g2_decap_8
XFILLER_42_170 VPWR VGND sg13g2_fill_1
X_2880_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\] net772 _0780_ _0390_
+ VPWR VGND sg13g2_mux2_1
X_4903__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_31_899 VPWR VGND sg13g2_decap_8
X_4550_ net680 net731 _0103_ VPWR VGND sg13g2_nor2_1
X_4481_ net670 net721 _0034_ VPWR VGND sg13g2_nor2_1
X_3501_ VGND VPWR _1229_ _1230_ _1231_ _1221_ sg13g2_a21oi_1
X_3432_ _1134_ VPWR _1162_ VGND _1145_ _1161_ sg13g2_o21ai_1
X_3363_ _1083_ _1092_ _1093_ VPWR VGND sg13g2_nor2_1
X_5102_ net797 VGND VPWR net695 serialize.n420\[6\] clknet_3_2__leaf_clk_regs sg13g2_dfrbpq_1
X_3294_ net611 videogen.fancy_shader.video_x\[3\] _1024_ VPWR VGND sg13g2_nor2_1
X_5033_ net279 VGND VPWR _0580_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\]
+ _0228_ sg13g2_dfrbpq_1
XFILLER_39_933 VPWR VGND sg13g2_decap_4
X_4984__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_41_608 VPWR VGND sg13g2_decap_4
XFILLER_15_38 VPWR VGND sg13g2_decap_4
XFILLER_34_682 VPWR VGND sg13g2_fill_2
X_4817_ net342 VGND VPWR _0368_ videogen.test_lut_thingy.gol_counter_reg\[2\] net643
+ sg13g2_dfrbpq_1
XFILLER_5_509 VPWR VGND sg13g2_fill_2
X_4748_ net95 VGND VPWR _0299_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\]
+ _0030_ sg13g2_dfrbpq_1
X_4679_ net686 net737 _0232_ VPWR VGND sg13g2_nor2_1
Xoutput15 net15 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_748 VPWR VGND sg13g2_decap_8
XFILLER_45_936 VPWR VGND sg13g2_decap_8
XFILLER_44_457 VPWR VGND sg13g2_decap_4
XFILLER_44_435 VPWR VGND sg13g2_fill_1
XFILLER_44_424 VPWR VGND sg13g2_decap_8
XFILLER_16_148 VPWR VGND sg13g2_fill_1
XFILLER_25_693 VPWR VGND sg13g2_decap_8
XFILLER_31_118 VPWR VGND sg13g2_fill_2
XFILLER_13_877 VPWR VGND sg13g2_decap_8
X_4820__339 VPWR VGND net339 sg13g2_tiehi
X_4939__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_9_848 VPWR VGND sg13g2_decap_8
XFILLER_9_859 VPWR VGND sg13g2_fill_2
XFILLER_13_888 VPWR VGND sg13g2_fill_1
X_4857__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_48_730 VPWR VGND sg13g2_fill_1
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_47_284 VPWR VGND sg13g2_fill_2
X_3981_ _1694_ _1697_ _1687_ _1707_ VPWR VGND sg13g2_nand3_1
X_2932_ videogen.fancy_shader.video_x\[8\] videogen.fancy_shader.video_x\[9\] _0791_
+ VPWR VGND sg13g2_and2_1
X_2863_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\] net761 _0777_ _0404_
+ VPWR VGND sg13g2_mux2_1
X_4602_ net666 net717 _0155_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
X_2794_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\] _0759_ _0455_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_195 VPWR VGND sg13g2_decap_8
XFILLER_8_870 VPWR VGND sg13g2_decap_8
X_4533_ net660 net711 _0086_ VPWR VGND sg13g2_nor2_1
X_4464_ net655 net706 _0017_ VPWR VGND sg13g2_nor2_1
X_4395_ _2084_ _2082_ _2086_ VPWR VGND sg13g2_xor2_1
X_3415_ VGND VPWR _1141_ _1143_ _1145_ _1056_ sg13g2_a21oi_1
X_3346_ _1076_ _1073_ _1075_ VPWR VGND sg13g2_xnor2_1
X_3277_ _1003_ VPWR _1007_ VGND _1004_ _1005_ sg13g2_o21ai_1
X_5016_ net94 VGND VPWR _0563_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\]
+ _0211_ sg13g2_dfrbpq_1
XFILLER_26_435 VPWR VGND sg13g2_fill_1
XFILLER_27_947 VPWR VGND sg13g2_decap_8
X_4726__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_41_449 VPWR VGND sg13g2_decap_8
XFILLER_35_991 VPWR VGND sg13g2_decap_8
XFILLER_22_652 VPWR VGND sg13g2_fill_1
XFILLER_10_814 VPWR VGND sg13g2_decap_8
XFILLER_10_847 VPWR VGND sg13g2_decap_8
X_4887__222 VPWR VGND net222 sg13g2_tiehi
XFILLER_29_273 VPWR VGND sg13g2_decap_8
XFILLER_29_284 VPWR VGND sg13g2_fill_2
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_41_972 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_8_122 VPWR VGND sg13g2_decap_4
XFILLER_9_667 VPWR VGND sg13g2_fill_2
XFILLER_32_80 VPWR VGND sg13g2_decap_4
X_4935__256 VPWR VGND net256 sg13g2_tiehi
X_3200_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] _0954_
+ _0956_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] sg13g2_a21oi_1
X_4180_ _1903_ _1901_ _1902_ VPWR VGND sg13g2_nand2b_1
X_3131_ _0909_ videogen.fancy_shader.video_x\[8\] _0906_ VPWR VGND sg13g2_xnor2_1
X_3062_ tmds_red.n100 tmds_red.n114 _0852_ VPWR VGND sg13g2_nor2_1
XFILLER_17_991 VPWR VGND sg13g2_decap_8
XFILLER_24_939 VPWR VGND sg13g2_decap_8
X_3964_ _1685_ _1689_ _1684_ _1690_ VPWR VGND sg13g2_nand3_1
XFILLER_23_449 VPWR VGND sg13g2_fill_2
X_2915_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\] net777 _0787_ _0288_
+ VPWR VGND sg13g2_mux2_1
X_3895_ _1251_ _1250_ _1621_ _0375_ VPWR VGND sg13g2_a21o_1
XFILLER_32_983 VPWR VGND sg13g2_decap_8
X_2846_ VPWR _0773_ _0772_ VGND sg13g2_inv_1
X_2777_ _0756_ _0702_ _0751_ VPWR VGND sg13g2_nand2_2
X_4516_ net674 net725 _0069_ VPWR VGND sg13g2_nor2_1
X_4447_ _2112_ _2134_ _2110_ _2136_ VPWR VGND sg13g2_nand3_1
Xfanout624 net625 net624 VPWR VGND sg13g2_buf_8
Xfanout613 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] net613 VPWR VGND
+ sg13g2_buf_8
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
Xfanout646 net649 net646 VPWR VGND sg13g2_buf_8
X_4378_ _0840_ _2071_ _2072_ VPWR VGND sg13g2_nor2_1
Xfanout657 net660 net657 VPWR VGND sg13g2_buf_8
Xfanout635 net639 net635 VPWR VGND sg13g2_buf_2
X_3329_ _1059_ _1043_ _1045_ VPWR VGND sg13g2_nand2_1
Xfanout679 net680 net679 VPWR VGND sg13g2_buf_8
Xfanout668 net673 net668 VPWR VGND sg13g2_buf_8
XFILLER_2_1014 VPWR VGND sg13g2_decap_8
XFILLER_39_582 VPWR VGND sg13g2_fill_1
XFILLER_27_722 VPWR VGND sg13g2_decap_4
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_26_243 VPWR VGND sg13g2_decap_4
XFILLER_27_788 VPWR VGND sg13g2_fill_1
XFILLER_30_909 VPWR VGND sg13g2_decap_8
XFILLER_23_983 VPWR VGND sg13g2_decap_8
XFILLER_6_626 VPWR VGND sg13g2_decap_8
XFILLER_6_604 VPWR VGND sg13g2_decap_4
XFILLER_2_832 VPWR VGND sg13g2_decap_8
XFILLER_49_324 VPWR VGND sg13g2_decap_8
XFILLER_18_722 VPWR VGND sg13g2_decap_4
XFILLER_18_766 VPWR VGND sg13g2_decap_4
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_14_950 VPWR VGND sg13g2_decap_8
X_2700_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\] _0739_ _0538_
+ VPWR VGND sg13g2_mux2_1
X_3680_ _1406_ _1407_ _1408_ _1409_ _1410_ VPWR VGND sg13g2_nor4_1
X_2631_ _0715_ _0720_ _0722_ VPWR VGND sg13g2_and2_1
X_2562_ VGND VPWR net592 _0674_ _0677_ net596 sg13g2_a21oi_1
X_4301_ _1991_ _1989_ _2002_ VPWR VGND sg13g2_nor2b_2
X_4232_ _1939_ _1929_ _1938_ VPWR VGND sg13g2_xnor2_1
X_4163_ _1872_ _1884_ _1886_ VPWR VGND sg13g2_and2_1
X_4094_ _1817_ _1112_ _1815_ VPWR VGND sg13g2_nand2b_1
X_3114_ _0899_ videogen.fancy_shader.video_x\[1\] net630 VPWR VGND sg13g2_xnor2_1
X_3045_ VGND VPWR net742 net434 _0265_ _0838_ sg13g2_a21oi_1
X_4996_ net211 VGND VPWR _0543_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\]
+ _0191_ sg13g2_dfrbpq_1
XFILLER_23_246 VPWR VGND sg13g2_decap_8
XFILLER_24_747 VPWR VGND sg13g2_decap_8
XFILLER_11_408 VPWR VGND sg13g2_decap_8
X_3947_ VPWR _1673_ _1672_ VGND sg13g2_inv_1
XFILLER_20_942 VPWR VGND sg13g2_decap_8
X_3878_ net593 VPWR _1607_ VGND _1605_ _1606_ sg13g2_o21ai_1
X_2829_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\] net783 _0768_ _0429_
+ VPWR VGND sg13g2_mux2_1
X_5014__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_3_607 VPWR VGND sg13g2_decap_8
XFILLER_2_139 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_48_68 VPWR VGND sg13g2_decap_8
XFILLER_46_316 VPWR VGND sg13g2_fill_2
XFILLER_46_327 VPWR VGND sg13g2_fill_2
XFILLER_27_552 VPWR VGND sg13g2_fill_2
XFILLER_42_533 VPWR VGND sg13g2_decap_4
XFILLER_42_566 VPWR VGND sg13g2_decap_8
XFILLER_30_717 VPWR VGND sg13g2_fill_2
XFILLER_11_942 VPWR VGND sg13g2_decap_8
XFILLER_23_791 VPWR VGND sg13g2_decap_8
XFILLER_7_968 VPWR VGND sg13g2_decap_8
XFILLER_10_463 VPWR VGND sg13g2_decap_8
X_4763__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_6_489 VPWR VGND sg13g2_decap_8
X_5032__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_1_194 VPWR VGND sg13g2_fill_2
XFILLER_46_872 VPWR VGND sg13g2_decap_8
X_4850_ net298 VGND VPWR _0401_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\]
+ _0058_ sg13g2_dfrbpq_1
XFILLER_33_533 VPWR VGND sg13g2_fill_2
X_3801_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\] net554 _1531_ VPWR
+ VGND sg13g2_nor2_1
X_4781_ net40 VGND VPWR _0332_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\]
+ net631 sg13g2_dfrbpq_2
X_3732_ net622 _1456_ _1461_ _1462_ VPWR VGND sg13g2_nor3_1
X_3663_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\] net561 _1393_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_294 VPWR VGND sg13g2_decap_8
X_2614_ _0680_ _0712_ _0713_ VPWR VGND sg13g2_nor2_2
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_3594_ net612 VPWR _1324_ VGND _1317_ _1323_ sg13g2_o21ai_1
X_2545_ videogen.fancy_shader.video_y\[8\] videogen.fancy_shader.video_y\[7\] _0632_
+ _0660_ VPWR VGND videogen.fancy_shader.video_y\[6\] sg13g2_nand4_1
X_4913__170 VPWR VGND net170 sg13g2_tiehi
X_4215_ net750 _1926_ _0498_ VPWR VGND sg13g2_nor2_1
X_4146_ _1867_ _1850_ _1851_ _1869_ VPWR VGND sg13g2_a21o_1
XFILLER_28_305 VPWR VGND sg13g2_decap_8
XFILLER_37_861 VPWR VGND sg13g2_fill_1
X_4077_ _1800_ _1726_ _1799_ VPWR VGND sg13g2_xnor2_1
X_3028_ net437 red_tmds_par\[3\] net697 serialize.n427\[3\] VPWR VGND sg13g2_mux2_1
XFILLER_36_393 VPWR VGND sg13g2_decap_8
XFILLER_34_48 VPWR VGND sg13g2_fill_1
X_4979_ net281 VGND VPWR _0526_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\]
+ _0174_ sg13g2_dfrbpq_1
XFILLER_24_599 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_3_3__leaf_clk_regs VGND sg13g2_inv_1
X_4966__355 VPWR VGND net355 sg13g2_tiehi
XFILLER_15_555 VPWR VGND sg13g2_fill_1
XFILLER_15_566 VPWR VGND sg13g2_fill_2
X_4973__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_6_231 VPWR VGND sg13g2_fill_1
X_4751__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_3_960 VPWR VGND sg13g2_decap_8
XFILLER_2_481 VPWR VGND sg13g2_decap_8
XFILLER_27_4 VPWR VGND sg13g2_fill_2
X_4000_ _1716_ VPWR _0378_ VGND _1722_ _1723_ sg13g2_o21ai_1
XFILLER_37_124 VPWR VGND sg13g2_fill_2
XFILLER_37_157 VPWR VGND sg13g2_decap_4
XFILLER_19_872 VPWR VGND sg13g2_decap_8
X_4902_ net192 VGND VPWR _0453_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\]
+ _0110_ sg13g2_dfrbpq_1
XFILLER_33_341 VPWR VGND sg13g2_fill_2
XFILLER_34_886 VPWR VGND sg13g2_decap_4
XFILLER_21_514 VPWR VGND sg13g2_decap_4
X_4833_ net326 VGND VPWR _0384_ red_tmds_par\[2\] net644 sg13g2_dfrbpq_1
X_4764_ net73 VGND VPWR _0315_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\]
+ _0036_ sg13g2_dfrbpq_1
X_3715_ net622 _1439_ _1444_ _1445_ VPWR VGND sg13g2_nor3_1
X_4695_ net662 net713 _0248_ VPWR VGND sg13g2_nor2_1
X_3646_ net614 VPWR _1376_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\]
+ net582 sg13g2_o21ai_1
X_3577_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\] net579 _1307_ VPWR
+ VGND sg13g2_nor2_1
X_2528_ VPWR _0646_ tmds_blue.dc_balancing_reg\[3\] VGND sg13g2_inv_1
Xhold37 serialize.n417\[7\] VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold15 serialize.n427\[6\] VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold26 serialize.n411\[2\] VPWR VGND net431 sg13g2_dlygate4sd3_1
X_4129_ VGND VPWR _1832_ _1836_ _1852_ _1835_ sg13g2_a21oi_1
XFILLER_29_658 VPWR VGND sg13g2_fill_1
XFILLER_45_14 VPWR VGND sg13g2_decap_4
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_16_308 VPWR VGND sg13g2_fill_1
XFILLER_40_878 VPWR VGND sg13g2_decap_4
XFILLER_20_580 VPWR VGND sg13g2_decap_8
XFILLER_10_94 VPWR VGND sg13g2_decap_4
XFILLER_48_923 VPWR VGND sg13g2_decap_8
XFILLER_47_400 VPWR VGND sg13g2_decap_8
XFILLER_0_996 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_decap_4
XFILLER_35_628 VPWR VGND sg13g2_fill_1
XFILLER_34_138 VPWR VGND sg13g2_decap_4
XFILLER_37_1025 VPWR VGND sg13g2_decap_4
X_4897__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_30_344 VPWR VGND sg13g2_decap_8
XFILLER_7_540 VPWR VGND sg13g2_fill_2
X_3500_ _1220_ _1225_ net545 _1230_ VPWR VGND sg13g2_nand3_1
X_4797__380 VPWR VGND net380 sg13g2_tiehi
XFILLER_30_399 VPWR VGND sg13g2_fill_1
X_4480_ net664 net715 _0033_ VPWR VGND sg13g2_nor2_1
XFILLER_7_573 VPWR VGND sg13g2_decap_8
XFILLER_7_562 VPWR VGND sg13g2_decap_8
X_3431_ VPWR VGND _1155_ _1147_ _1153_ _1032_ _1161_ _1033_ sg13g2_a221oi_1
X_3362_ _1092_ _1091_ _1090_ VPWR VGND sg13g2_nand2b_1
X_5101_ net800 VGND VPWR net416 serialize.n420\[4\] clknet_3_3__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_39_912 VPWR VGND sg13g2_fill_1
X_3293_ _1023_ net611 videogen.fancy_shader.video_x\[3\] VPWR VGND sg13g2_nand2_1
X_5032_ net287 VGND VPWR _0579_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\]
+ _0227_ sg13g2_dfrbpq_1
XFILLER_38_466 VPWR VGND sg13g2_fill_1
XFILLER_40_108 VPWR VGND sg13g2_fill_2
XFILLER_22_845 VPWR VGND sg13g2_fill_1
X_4816_ net343 VGND VPWR _0367_ videogen.test_lut_thingy.gol_counter_reg\[1\] net643
+ sg13g2_dfrbpq_2
XFILLER_21_366 VPWR VGND sg13g2_fill_1
X_4747_ net97 VGND VPWR _0298_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\]
+ _0029_ sg13g2_dfrbpq_1
X_4678_ net672 net722 _0231_ VPWR VGND sg13g2_nor2_1
X_3629_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\] net579 _1359_ VPWR
+ VGND sg13g2_nor2_1
Xoutput16 net16 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_727 VPWR VGND sg13g2_decap_8
XFILLER_0_226 VPWR VGND sg13g2_fill_1
XFILLER_5_1023 VPWR VGND sg13g2_decap_4
XFILLER_45_915 VPWR VGND sg13g2_decap_8
XFILLER_44_403 VPWR VGND sg13g2_decap_4
XFILLER_13_823 VPWR VGND sg13g2_fill_1
XFILLER_24_171 VPWR VGND sg13g2_fill_2
XFILLER_12_333 VPWR VGND sg13g2_decap_4
XFILLER_4_565 VPWR VGND sg13g2_decap_8
XFILLER_21_93 VPWR VGND sg13g2_fill_1
XFILLER_0_793 VPWR VGND sg13g2_decap_8
X_3980_ _1702_ _1705_ _1706_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_469 VPWR VGND sg13g2_decap_8
XFILLER_44_981 VPWR VGND sg13g2_decap_8
X_2931_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\] _0790_ _0267_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_160 VPWR VGND sg13g2_decap_4
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_2862_ _0721_ _0725_ _0777_ VPWR VGND sg13g2_nor2_2
X_4601_ net663 net714 _0154_ VPWR VGND sg13g2_nor2_1
XFILLER_31_675 VPWR VGND sg13g2_fill_1
X_2793_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\] _0759_ _0456_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_174 VPWR VGND sg13g2_decap_8
X_4532_ net657 net708 _0085_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_4719__145 VPWR VGND net145 sg13g2_tiehi
X_4463_ net668 net720 _0016_ VPWR VGND sg13g2_nor2_1
X_3414_ VPWR _1144_ _1143_ VGND sg13g2_inv_1
X_4394_ _2082_ _2084_ _2085_ VPWR VGND sg13g2_nor2_1
X_3345_ _1075_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.video_x\[6\]
+ VPWR VGND sg13g2_xnor2_1
X_3276_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_y\[1\] _1006_
+ VPWR VGND sg13g2_xor2_1
X_5015_ net102 VGND VPWR _0562_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\]
+ _0210_ sg13g2_dfrbpq_1
XFILLER_27_926 VPWR VGND sg13g2_decap_8
XFILLER_35_970 VPWR VGND sg13g2_fill_2
X_5023__381 VPWR VGND net381 sg13g2_tiehi
XFILLER_21_130 VPWR VGND sg13g2_fill_1
XFILLER_22_675 VPWR VGND sg13g2_decap_8
XFILLER_6_819 VPWR VGND sg13g2_decap_8
XFILLER_5_329 VPWR VGND sg13g2_fill_1
XFILLER_27_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_18_959 VPWR VGND sg13g2_decap_8
X_4924__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_32_417 VPWR VGND sg13g2_fill_1
XFILLER_41_951 VPWR VGND sg13g2_decap_8
XFILLER_41_940 VPWR VGND sg13g2_fill_2
XFILLER_13_642 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_145 VPWR VGND sg13g2_decap_8
XFILLER_8_156 VPWR VGND sg13g2_fill_1
X_3130_ _0908_ videogen.fancy_shader.video_x\[8\] _0906_ VPWR VGND sg13g2_nand2_1
XFILLER_0_590 VPWR VGND sg13g2_fill_2
X_3061_ tmds_red.n126 tmds_red.n132 _0851_ VPWR VGND sg13g2_nor2_1
XFILLER_48_583 VPWR VGND sg13g2_decap_8
XFILLER_35_222 VPWR VGND sg13g2_decap_4
XFILLER_24_918 VPWR VGND sg13g2_decap_8
XFILLER_17_970 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_4
XFILLER_35_288 VPWR VGND sg13g2_fill_2
X_3963_ _1675_ _1687_ _1689_ VPWR VGND sg13g2_nor2_1
X_4803__368 VPWR VGND net368 sg13g2_tiehi
X_2914_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\] net768 _0787_ _0289_
+ VPWR VGND sg13g2_mux2_1
X_3894_ _1549_ _1620_ _1621_ VPWR VGND sg13g2_and2_1
XFILLER_32_962 VPWR VGND sg13g2_decap_8
X_2845_ _0772_ _0680_ _0761_ VPWR VGND sg13g2_nand2_2
X_4515_ net675 net725 _0068_ VPWR VGND sg13g2_nor2_1
X_2776_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\] _0755_ _0469_
+ VPWR VGND sg13g2_mux2_1
X_4446_ VGND VPWR _2110_ _2112_ _2135_ _2134_ sg13g2_a21oi_1
X_4377_ VGND VPWR _2065_ _2070_ _2071_ _0847_ sg13g2_a21oi_1
Xfanout614 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net614 VPWR VGND
+ sg13g2_buf_8
Xfanout603 tmds_green.n100 net603 VPWR VGND sg13g2_buf_2
X_3328_ videogen.fancy_shader.video_x\[5\] videogen.fancy_shader.n646\[5\] _1058_
+ VPWR VGND sg13g2_xor2_1
Xfanout625 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\] net625 VPWR VGND
+ sg13g2_buf_8
Xfanout658 net660 net658 VPWR VGND sg13g2_buf_1
Xfanout636 net639 net636 VPWR VGND sg13g2_buf_8
Xfanout647 net649 net647 VPWR VGND sg13g2_buf_8
Xfanout669 net673 net669 VPWR VGND sg13g2_buf_2
X_3259_ VGND VPWR videogen.fancy_shader.video_y\[9\] _0993_ _0995_ _0981_ sg13g2_a21oi_1
XFILLER_26_288 VPWR VGND sg13g2_fill_2
XFILLER_41_236 VPWR VGND sg13g2_decap_4
XFILLER_14_439 VPWR VGND sg13g2_decap_4
XFILLER_23_962 VPWR VGND sg13g2_decap_8
XFILLER_5_115 VPWR VGND sg13g2_decap_8
X_4969__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_49_303 VPWR VGND sg13g2_decap_8
XFILLER_2_888 VPWR VGND sg13g2_decap_8
XFILLER_1_354 VPWR VGND sg13g2_fill_2
XFILLER_45_542 VPWR VGND sg13g2_fill_1
XFILLER_17_244 VPWR VGND sg13g2_fill_2
XFILLER_17_277 VPWR VGND sg13g2_fill_2
XFILLER_13_483 VPWR VGND sg13g2_fill_2
X_2630_ VGND VPWR _0721_ _0687_ _0680_ sg13g2_or2_1
XFILLER_9_498 VPWR VGND sg13g2_decap_8
X_2561_ net614 net619 net583 _0676_ VPWR VGND sg13g2_nor3_2
X_4300_ _2001_ tmds_blue.n126 _1996_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_181 VPWR VGND sg13g2_decap_8
X_4231_ _1938_ _1932_ _1936_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_74 VPWR VGND sg13g2_fill_1
X_4162_ _1872_ _1884_ _1885_ VPWR VGND sg13g2_nor2_1
X_4093_ _1816_ net542 _1815_ VPWR VGND sg13g2_nand2_1
X_3113_ net630 _0898_ _0303_ VPWR VGND sg13g2_nor2_1
XFILLER_28_509 VPWR VGND sg13g2_decap_8
X_3044_ net794 VPWR _0838_ VGND net741 net434 sg13g2_o21ai_1
XFILLER_24_726 VPWR VGND sg13g2_decap_8
X_4995_ net215 VGND VPWR _0542_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\]
+ _0190_ sg13g2_dfrbpq_1
XFILLER_23_236 VPWR VGND sg13g2_fill_1
X_3946_ _1660_ VPWR _1672_ VGND _1666_ _1669_ sg13g2_o21ai_1
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
XFILLER_20_921 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_fill_2
X_3877_ _1562_ VPWR _1606_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\]
+ net551 sg13g2_o21ai_1
X_2828_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\] net773 _0768_ _0430_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_998 VPWR VGND sg13g2_decap_8
X_2759_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\] _0752_ _0483_
+ VPWR VGND sg13g2_mux2_1
X_4429_ _2118_ _2114_ _2119_ VPWR VGND sg13g2_xor2_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1016 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_339 VPWR VGND sg13g2_fill_2
XFILLER_39_391 VPWR VGND sg13g2_decap_8
XFILLER_27_542 VPWR VGND sg13g2_decap_4
XFILLER_42_512 VPWR VGND sg13g2_fill_2
XFILLER_15_715 VPWR VGND sg13g2_decap_4
XFILLER_27_586 VPWR VGND sg13g2_decap_8
XFILLER_11_921 VPWR VGND sg13g2_decap_8
XFILLER_6_402 VPWR VGND sg13g2_decap_8
XFILLER_7_947 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
X_4748__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_2_641 VPWR VGND sg13g2_fill_1
XFILLER_2_652 VPWR VGND sg13g2_fill_1
XFILLER_49_155 VPWR VGND sg13g2_fill_1
XFILLER_38_829 VPWR VGND sg13g2_fill_2
XFILLER_49_188 VPWR VGND sg13g2_decap_8
XFILLER_46_851 VPWR VGND sg13g2_decap_4
X_4780_ net42 VGND VPWR _0331_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\]
+ net632 sg13g2_dfrbpq_2
X_3800_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\] net563 _1530_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_21_718 VPWR VGND sg13g2_decap_8
X_4722__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_20_239 VPWR VGND sg13g2_decap_8
X_3731_ _1457_ _1458_ _1459_ _1460_ _1461_ VPWR VGND sg13g2_nor4_1
X_3662_ net596 VPWR _1392_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\]
+ net574 sg13g2_o21ai_1
X_3593_ net615 VPWR _1323_ VGND _1318_ _1322_ sg13g2_o21ai_1
X_2613_ _0712_ _0686_ VPWR VGND _0682_ sg13g2_nand2b_2
X_2544_ _0659_ VPWR _0262_ VGND net444 serialize.n433\[1\] sg13g2_o21ai_1
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_4214_ VGND VPWR _0844_ _0848_ _1926_ _1925_ sg13g2_a21oi_1
X_4145_ VGND VPWR _1850_ _1867_ _1868_ _1851_ sg13g2_a21oi_1
X_5077__47 VPWR VGND net47 sg13g2_tiehi
X_4076_ _1031_ _1797_ _1799_ VPWR VGND sg13g2_and2_1
XFILLER_37_884 VPWR VGND sg13g2_decap_8
X_3027_ net431 red_tmds_par\[2\] net697 serialize.n427\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_36_350 VPWR VGND sg13g2_fill_2
XFILLER_24_567 VPWR VGND sg13g2_decap_4
X_4978_ net285 VGND VPWR _0525_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\]
+ _0173_ sg13g2_dfrbpq_1
X_3929_ _1637_ _1644_ _1655_ VPWR VGND sg13g2_nor2_1
Xclkload4 clknet_3_4__leaf_clk_regs clkload4/X VPWR VGND sg13g2_buf_1
XFILLER_20_762 VPWR VGND sg13g2_decap_4
X_4760__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
XFILLER_47_604 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_fill_2
XFILLER_43_832 VPWR VGND sg13g2_decap_8
XFILLER_42_331 VPWR VGND sg13g2_decap_4
XFILLER_27_394 VPWR VGND sg13g2_fill_1
XFILLER_42_386 VPWR VGND sg13g2_fill_2
XFILLER_30_526 VPWR VGND sg13g2_decap_8
XFILLER_11_751 VPWR VGND sg13g2_decap_8
XFILLER_11_762 VPWR VGND sg13g2_fill_2
XFILLER_10_294 VPWR VGND sg13g2_decap_8
XFILLER_7_788 VPWR VGND sg13g2_decap_8
XFILLER_2_471 VPWR VGND sg13g2_fill_2
XFILLER_38_615 VPWR VGND sg13g2_decap_8
X_4867__265 VPWR VGND net265 sg13g2_tiehi
XFILLER_19_840 VPWR VGND sg13g2_decap_8
XFILLER_18_394 VPWR VGND sg13g2_fill_1
X_4901_ net194 VGND VPWR _0452_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[3\]
+ _0109_ sg13g2_dfrbpq_1
XFILLER_33_320 VPWR VGND sg13g2_decap_8
XFILLER_34_865 VPWR VGND sg13g2_decap_8
XFILLER_21_537 VPWR VGND sg13g2_fill_1
X_4832_ net327 VGND VPWR _0383_ tmds_red.n132 net640 sg13g2_dfrbpq_2
XFILLER_34_898 VPWR VGND sg13g2_fill_2
X_4763_ net75 VGND VPWR _0314_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\]
+ _0035_ sg13g2_dfrbpq_1
X_4694_ net665 net716 _0247_ VPWR VGND sg13g2_nor2_1
X_3714_ _1440_ _1441_ _1442_ _1443_ _1444_ VPWR VGND sg13g2_nor4_1
X_4874__247 VPWR VGND net247 sg13g2_tiehi
X_3645_ _1375_ net613 _1374_ VPWR VGND sg13g2_nand2b_1
X_3576_ _1302_ _1303_ _1304_ _1305_ _1306_ VPWR VGND sg13g2_nor4_1
XFILLER_1_909 VPWR VGND sg13g2_decap_8
X_2527_ VPWR _0645_ tmds_blue.dc_balancing_reg\[1\] VGND sg13g2_inv_1
Xhold16 serialize.n414\[5\] VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold38 serialize.n417\[4\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold27 serialize.n411\[1\] VPWR VGND net432 sg13g2_dlygate4sd3_1
XFILLER_29_38 VPWR VGND sg13g2_fill_2
XFILLER_29_604 VPWR VGND sg13g2_fill_2
X_4846__305 VPWR VGND net305 sg13g2_tiehi
X_4128_ _1851_ _1848_ _1849_ _1844_ _1839_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_147 VPWR VGND sg13g2_decap_4
XFILLER_45_26 VPWR VGND sg13g2_fill_2
X_4059_ _1782_ _1774_ _1781_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_386 VPWR VGND sg13g2_decap_8
XFILLER_4_736 VPWR VGND sg13g2_decap_4
XFILLER_10_51 VPWR VGND sg13g2_decap_8
Xclkbuf_regs_0_clk clk clk_regs VPWR VGND sg13g2_buf_8
XFILLER_3_279 VPWR VGND sg13g2_fill_1
XFILLER_48_902 VPWR VGND sg13g2_decap_8
XFILLER_0_975 VPWR VGND sg13g2_decap_8
XFILLER_48_979 VPWR VGND sg13g2_decap_8
XFILLER_19_147 VPWR VGND sg13g2_fill_2
XFILLER_47_489 VPWR VGND sg13g2_decap_4
XFILLER_19_169 VPWR VGND sg13g2_fill_1
XFILLER_35_618 VPWR VGND sg13g2_fill_2
XFILLER_16_843 VPWR VGND sg13g2_decap_8
XFILLER_28_692 VPWR VGND sg13g2_decap_8
XFILLER_37_1004 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_fill_2
XFILLER_43_684 VPWR VGND sg13g2_decap_8
XFILLER_43_673 VPWR VGND sg13g2_decap_8
XFILLER_42_194 VPWR VGND sg13g2_decap_4
XFILLER_15_397 VPWR VGND sg13g2_decap_8
XFILLER_30_367 VPWR VGND sg13g2_fill_1
X_3430_ _1157_ _1159_ _1160_ VPWR VGND _1156_ sg13g2_nand3b_1
X_3361_ VGND VPWR _1091_ videogen.fancy_shader.n646\[7\] videogen.fancy_shader.video_y\[7\]
+ sg13g2_or2_1
X_5100_ net800 VGND VPWR serialize.n431\[5\] serialize.n420\[3\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_791 VPWR VGND sg13g2_decap_8
X_5031_ net295 VGND VPWR _0578_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\]
+ _0226_ sg13g2_dfrbpq_1
X_3292_ VPWR _1022_ net545 VGND sg13g2_inv_1
XFILLER_39_979 VPWR VGND sg13g2_decap_8
XFILLER_38_478 VPWR VGND sg13g2_decap_8
XFILLER_25_106 VPWR VGND sg13g2_fill_2
XFILLER_26_629 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_fill_2
XFILLER_22_824 VPWR VGND sg13g2_decap_8
XFILLER_34_684 VPWR VGND sg13g2_fill_1
XFILLER_21_345 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
X_4815_ net344 VGND VPWR _0366_ videogen.test_lut_thingy.gol_counter_reg\[0\] net643
+ sg13g2_dfrbpq_2
X_5056__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_21_356 VPWR VGND sg13g2_fill_2
XFILLER_21_378 VPWR VGND sg13g2_decap_4
X_4746_ net99 VGND VPWR _0297_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\]
+ _0028_ sg13g2_dfrbpq_1
X_4677_ net671 net722 _0230_ VPWR VGND sg13g2_nor2_1
X_3628_ net598 VPWR _1358_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\]
+ net555 sg13g2_o21ai_1
Xoutput17 net17 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_706 VPWR VGND sg13g2_decap_8
X_3559_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\] net566 _1289_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_205 VPWR VGND sg13g2_decap_8
X_4813__348 VPWR VGND net348 sg13g2_tiehi
XFILLER_0_249 VPWR VGND sg13g2_decap_8
XFILLER_5_1002 VPWR VGND sg13g2_decap_8
XFILLER_17_607 VPWR VGND sg13g2_fill_2
XFILLER_17_629 VPWR VGND sg13g2_fill_2
XFILLER_24_183 VPWR VGND sg13g2_fill_1
XFILLER_9_828 VPWR VGND sg13g2_decap_4
XFILLER_12_356 VPWR VGND sg13g2_decap_8
XFILLER_40_698 VPWR VGND sg13g2_decap_4
XFILLER_21_61 VPWR VGND sg13g2_fill_1
XFILLER_0_772 VPWR VGND sg13g2_decap_8
XFILLER_48_754 VPWR VGND sg13g2_fill_2
XFILLER_47_231 VPWR VGND sg13g2_fill_1
XFILLER_36_938 VPWR VGND sg13g2_fill_2
XFILLER_47_286 VPWR VGND sg13g2_fill_1
XFILLER_44_960 VPWR VGND sg13g2_decap_8
X_2930_ net778 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\] _0790_ _0268_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_673 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_fill_1
XFILLER_31_621 VPWR VGND sg13g2_decap_8
X_2861_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\] net787 _0776_ _0405_
+ VPWR VGND sg13g2_mux2_1
X_4600_ net654 net705 _0153_ VPWR VGND sg13g2_nor2_1
X_2792_ _0759_ _0727_ _0751_ VPWR VGND sg13g2_nand2_2
XFILLER_30_186 VPWR VGND sg13g2_fill_1
X_4531_ net657 net708 _0084_ VPWR VGND sg13g2_nor2_1
X_4462_ net659 net710 _0015_ VPWR VGND sg13g2_nor2_1
X_3413_ _1130_ _1128_ _1142_ _1143_ VPWR VGND sg13g2_a21o_1
X_4393_ _2083_ VPWR _2084_ VGND tmds_blue.dc_balancing_reg\[1\] _2076_ sg13g2_o21ai_1
X_3344_ _1074_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.video_x\[6\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3275_ net608 videogen.fancy_shader.n646\[1\] _1005_ VPWR VGND sg13g2_nor2_1
X_5014_ net110 VGND VPWR _0561_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\]
+ _0209_ sg13g2_dfrbpq_1
XFILLER_38_264 VPWR VGND sg13g2_fill_1
XFILLER_38_231 VPWR VGND sg13g2_decap_4
XFILLER_27_905 VPWR VGND sg13g2_decap_8
XFILLER_41_429 VPWR VGND sg13g2_fill_2
X_4729_ net133 VGND VPWR _0280_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[1\]
+ _0011_ sg13g2_dfrbpq_1
XFILLER_27_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
XFILLER_44_212 VPWR VGND sg13g2_fill_2
XFILLER_17_437 VPWR VGND sg13g2_fill_2
XFILLER_18_938 VPWR VGND sg13g2_decap_8
XFILLER_33_908 VPWR VGND sg13g2_fill_2
XFILLER_26_982 VPWR VGND sg13g2_decap_8
XFILLER_25_492 VPWR VGND sg13g2_fill_1
XFILLER_34_1007 VPWR VGND sg13g2_decap_8
X_5035__264 VPWR VGND net264 sg13g2_tiehi
XFILLER_5_853 VPWR VGND sg13g2_decap_8
XFILLER_5_897 VPWR VGND sg13g2_decap_8
X_3060_ VGND VPWR tmds_red.n126 tmds_red.n132 _0850_ tmds_red.n102 sg13g2_a21oi_1
XFILLER_48_562 VPWR VGND sg13g2_decap_8
XFILLER_16_470 VPWR VGND sg13g2_fill_1
X_3962_ _1623_ _1021_ _1688_ VPWR VGND sg13g2_xor2_1
XFILLER_32_930 VPWR VGND sg13g2_decap_8
X_2913_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\] net756 _0787_ _0290_
+ VPWR VGND sg13g2_mux2_1
X_3893_ _1449_ _1616_ _1352_ _1620_ VPWR VGND sg13g2_nand3_1
X_2844_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\] net783 _0771_ _0417_
+ VPWR VGND sg13g2_mux2_1
X_4514_ net674 net727 _0067_ VPWR VGND sg13g2_nor2_1
X_2775_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\] _0755_ _0470_
+ VPWR VGND sg13g2_mux2_1
X_4445_ _2134_ tmds_blue.dc_balancing_reg\[4\] _2133_ VPWR VGND sg13g2_xnor2_1
X_4376_ _2070_ _2067_ _2069_ VPWR VGND sg13g2_xnor2_1
Xfanout615 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net615 VPWR VGND
+ sg13g2_buf_8
Xfanout604 net605 net604 VPWR VGND sg13g2_buf_8
Xfanout648 net649 net648 VPWR VGND sg13g2_buf_1
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_8
X_3327_ _1057_ _0634_ _0640_ VPWR VGND sg13g2_nand2_1
Xfanout637 net639 net637 VPWR VGND sg13g2_buf_2
Xfanout659 net660 net659 VPWR VGND sg13g2_buf_8
X_3258_ videogen.fancy_shader.video_y\[9\] _0993_ _0994_ VPWR VGND sg13g2_nor2_1
X_3189_ _0944_ _0949_ _0332_ VPWR VGND sg13g2_nor2_1
XFILLER_23_941 VPWR VGND sg13g2_decap_8
XFILLER_10_602 VPWR VGND sg13g2_decap_8
X_4775__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_10_646 VPWR VGND sg13g2_decap_8
XFILLER_2_801 VPWR VGND sg13g2_decap_8
XFILLER_2_867 VPWR VGND sg13g2_decap_8
XFILLER_49_359 VPWR VGND sg13g2_decap_8
XFILLER_32_237 VPWR VGND sg13g2_decap_8
XFILLER_41_760 VPWR VGND sg13g2_decap_4
XFILLER_14_985 VPWR VGND sg13g2_decap_8
XFILLER_43_70 VPWR VGND sg13g2_fill_1
X_2560_ VGND VPWR _0675_ net626 net624 sg13g2_or2_1
XFILLER_5_672 VPWR VGND sg13g2_decap_8
XFILLER_4_160 VPWR VGND sg13g2_fill_2
XFILLER_4_31 VPWR VGND sg13g2_decap_8
X_4230_ _1932_ _1936_ _1937_ VPWR VGND sg13g2_nor2b_1
X_4161_ _1875_ _1883_ _1884_ VPWR VGND sg13g2_nor2b_1
X_4092_ _1810_ _1738_ _1815_ VPWR VGND sg13g2_xor2_1
X_3112_ _0898_ net795 VPWR VGND _0897_ sg13g2_nand2b_2
X_3043_ tmds_blue.dc_balancing_reg\[0\] _0836_ _0264_ VPWR VGND sg13g2_and2_1
X_4994_ net219 VGND VPWR _0541_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\]
+ _0189_ sg13g2_dfrbpq_1
X_3945_ VGND VPWR _1671_ _1670_ _1666_ sg13g2_or2_1
XFILLER_23_18 VPWR VGND sg13g2_fill_2
XFILLER_20_977 VPWR VGND sg13g2_decap_8
X_3876_ _1563_ VPWR _1605_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\]
+ net573 sg13g2_o21ai_1
X_2827_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\] net768 _0768_ _0431_
+ VPWR VGND sg13g2_mux2_1
X_2758_ net756 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\] _0752_ _0484_
+ VPWR VGND sg13g2_mux2_1
X_4428_ _2118_ _2116_ _2117_ VPWR VGND sg13g2_nand2_1
X_2689_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\] _0737_ _0547_
+ VPWR VGND sg13g2_mux2_1
X_4359_ _2054_ _2051_ _2053_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_318 VPWR VGND sg13g2_fill_1
XFILLER_39_370 VPWR VGND sg13g2_decap_4
XFILLER_27_565 VPWR VGND sg13g2_decap_8
XFILLER_14_226 VPWR VGND sg13g2_decap_8
XFILLER_14_248 VPWR VGND sg13g2_decap_8
XFILLER_30_719 VPWR VGND sg13g2_fill_1
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_22_281 VPWR VGND sg13g2_decap_8
XFILLER_10_454 VPWR VGND sg13g2_decap_4
XFILLER_10_476 VPWR VGND sg13g2_fill_1
XFILLER_10_487 VPWR VGND sg13g2_fill_2
XFILLER_6_458 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_1_174 VPWR VGND sg13g2_fill_1
XFILLER_49_134 VPWR VGND sg13g2_decap_8
XFILLER_49_167 VPWR VGND sg13g2_decap_8
XFILLER_18_565 VPWR VGND sg13g2_fill_1
XFILLER_45_395 VPWR VGND sg13g2_fill_2
XFILLER_45_373 VPWR VGND sg13g2_fill_2
XFILLER_14_793 VPWR VGND sg13g2_decap_8
X_3730_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\] net589 _1460_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_13_281 VPWR VGND sg13g2_decap_8
X_3661_ _1387_ _1388_ _1389_ _1390_ _1391_ VPWR VGND sg13g2_nor4_1
X_3592_ _1321_ VPWR _1322_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\]
+ net551 sg13g2_o21ai_1
X_2612_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\] _0711_ _0598_
+ VPWR VGND sg13g2_mux2_1
X_2543_ _0659_ net444 _0658_ VPWR VGND sg13g2_nand2_1
XFILLER_6_970 VPWR VGND sg13g2_decap_8
X_4213_ net607 VPWR _1925_ VGND tmds_green.n126 _0844_ sg13g2_o21ai_1
X_4144_ _1845_ VPWR _1867_ VGND _1851_ _1853_ sg13g2_o21ai_1
X_4075_ _1798_ _1021_ _1796_ VPWR VGND sg13g2_xnor2_1
X_3026_ net432 red_tmds_par\[1\] net698 serialize.n427\[1\] VPWR VGND sg13g2_mux2_1
XFILLER_24_513 VPWR VGND sg13g2_fill_2
XFILLER_34_17 VPWR VGND sg13g2_fill_1
XFILLER_34_28 VPWR VGND sg13g2_fill_2
XFILLER_12_719 VPWR VGND sg13g2_decap_4
X_4977_ net289 VGND VPWR _0524_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\]
+ _0172_ sg13g2_dfrbpq_1
Xclkload5 VPWR clkload5/Y clknet_3_5__leaf_clk_regs VGND sg13g2_inv_1
X_3928_ _1635_ _1643_ _1647_ _1649_ _1654_ VPWR VGND sg13g2_or4_1
XFILLER_32_590 VPWR VGND sg13g2_fill_2
X_3859_ _1586_ VPWR _1588_ VGND net621 _1587_ sg13g2_o21ai_1
XFILLER_30_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_929 VPWR VGND sg13g2_decap_8
XFILLER_28_852 VPWR VGND sg13g2_fill_2
XFILLER_42_354 VPWR VGND sg13g2_fill_1
XFILLER_15_546 VPWR VGND sg13g2_fill_2
X_4999__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_30_505 VPWR VGND sg13g2_decap_8
XFILLER_11_730 VPWR VGND sg13g2_fill_1
XFILLER_23_590 VPWR VGND sg13g2_decap_8
XFILLER_7_723 VPWR VGND sg13g2_decap_4
XFILLER_11_785 VPWR VGND sg13g2_decap_8
XFILLER_6_255 VPWR VGND sg13g2_decap_8
XFILLER_3_995 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_27_6 VPWR VGND sg13g2_fill_1
XFILLER_18_351 VPWR VGND sg13g2_decap_8
XFILLER_45_170 VPWR VGND sg13g2_fill_2
X_4900_ net196 VGND VPWR _0451_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\]
+ _0108_ sg13g2_dfrbpq_1
XFILLER_18_384 VPWR VGND sg13g2_decap_4
XFILLER_34_844 VPWR VGND sg13g2_decap_8
X_4831_ net328 VGND VPWR _0382_ tmds_red.n126 net644 sg13g2_dfrbpq_2
X_5039__229 VPWR VGND net229 sg13g2_tiehi
XFILLER_33_387 VPWR VGND sg13g2_decap_4
X_4762_ net77 VGND VPWR _0313_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\]
+ _0034_ sg13g2_dfrbpq_1
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_4693_ net661 net712 _0246_ VPWR VGND sg13g2_nor2_1
X_3713_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\] net580 _1443_ VPWR
+ VGND sg13g2_nor2_1
X_3644_ net592 _1368_ _1373_ _1374_ VPWR VGND sg13g2_nor3_1
X_3575_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\] net579 _1305_ VPWR
+ VGND sg13g2_nor2_1
X_2526_ VPWR _0644_ tmds_blue.dc_balancing_reg\[4\] VGND sg13g2_inv_1
X_4750__91 VPWR VGND net91 sg13g2_tiehi
Xhold28 serialize.n417\[0\] VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold17 serialize.n414\[4\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold39 _0004_ VPWR VGND net444 sg13g2_dlygate4sd3_1
X_4127_ _1848_ _1849_ _1850_ VPWR VGND sg13g2_and2_1
XFILLER_37_660 VPWR VGND sg13g2_decap_8
X_4058_ _1781_ _1762_ _1767_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_800 VPWR VGND sg13g2_fill_2
X_5061__260 VPWR VGND net260 sg13g2_tiehi
X_3009_ net445 blue_tmds_par\[5\] net695 serialize.n429\[5\] VPWR VGND sg13g2_mux2_1
XFILLER_24_321 VPWR VGND sg13g2_fill_2
XFILLER_25_899 VPWR VGND sg13g2_decap_8
XFILLER_12_538 VPWR VGND sg13g2_fill_1
XFILLER_4_715 VPWR VGND sg13g2_decap_8
X_4736__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_10_30 VPWR VGND sg13g2_decap_8
XFILLER_0_954 VPWR VGND sg13g2_decap_8
X_4927__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_48_958 VPWR VGND sg13g2_decap_8
XFILLER_47_446 VPWR VGND sg13g2_fill_2
XFILLER_16_800 VPWR VGND sg13g2_fill_2
XFILLER_34_107 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_fill_2
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_27_192 VPWR VGND sg13g2_decap_4
XFILLER_16_888 VPWR VGND sg13g2_fill_2
XFILLER_31_825 VPWR VGND sg13g2_decap_8
XFILLER_7_597 VPWR VGND sg13g2_fill_1
X_3360_ videogen.fancy_shader.video_y\[7\] videogen.fancy_shader.n646\[7\] _1090_
+ VPWR VGND sg13g2_and2_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
XFILLER_3_770 VPWR VGND sg13g2_fill_1
X_5030_ net302 VGND VPWR _0577_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\]
+ _0225_ sg13g2_dfrbpq_1
X_3291_ _1019_ _1020_ _1021_ VPWR VGND sg13g2_and2_1
XFILLER_19_682 VPWR VGND sg13g2_fill_1
XFILLER_15_19 VPWR VGND sg13g2_fill_2
XFILLER_22_803 VPWR VGND sg13g2_decap_8
XFILLER_33_162 VPWR VGND sg13g2_decap_8
XFILLER_34_696 VPWR VGND sg13g2_decap_8
X_4814_ net346 VGND VPWR _0365_ videogen.fancy_shader.video_y\[9\] net635 sg13g2_dfrbpq_2
XFILLER_21_313 VPWR VGND sg13g2_fill_1
X_4745_ net101 VGND VPWR _0296_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\]
+ _0027_ sg13g2_dfrbpq_1
X_4676_ net671 net722 _0229_ VPWR VGND sg13g2_nor2_1
X_4956__389 VPWR VGND net389 sg13g2_tiehi
X_3627_ _1353_ _1354_ _1355_ _1356_ _1357_ VPWR VGND sg13g2_nor4_1
X_3558_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\] net589 _1288_ VPWR
+ VGND sg13g2_nor2_1
Xoutput18 net18 uo_out[5] VPWR VGND sg13g2_buf_1
X_3489_ VGND VPWR _1219_ _1218_ _1217_ sg13g2_or2_1
XFILLER_29_402 VPWR VGND sg13g2_decap_8
XFILLER_40_622 VPWR VGND sg13g2_fill_1
XFILLER_13_847 VPWR VGND sg13g2_decap_4
XFILLER_24_195 VPWR VGND sg13g2_decap_8
XFILLER_12_379 VPWR VGND sg13g2_fill_2
XFILLER_21_891 VPWR VGND sg13g2_decap_8
XFILLER_4_545 VPWR VGND sg13g2_fill_2
XFILLER_0_751 VPWR VGND sg13g2_decap_8
XFILLER_36_928 VPWR VGND sg13g2_fill_1
XFILLER_35_427 VPWR VGND sg13g2_fill_1
XFILLER_35_438 VPWR VGND sg13g2_decap_8
XFILLER_43_493 VPWR VGND sg13g2_fill_1
X_2860_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\] net777 _0776_ _0406_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_184 VPWR VGND sg13g2_decap_8
XFILLER_31_644 VPWR VGND sg13g2_fill_2
XFILLER_30_143 VPWR VGND sg13g2_decap_4
XFILLER_12_880 VPWR VGND sg13g2_decap_8
X_2791_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\] net788 _0758_ _0457_
+ VPWR VGND sg13g2_mux2_1
X_4530_ net657 net708 _0083_ VPWR VGND sg13g2_nor2_1
XFILLER_11_390 VPWR VGND sg13g2_decap_4
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_7_372 VPWR VGND sg13g2_decap_4
XFILLER_7_75 VPWR VGND sg13g2_decap_8
X_4461_ net663 net714 _0014_ VPWR VGND sg13g2_nor2_1
X_3412_ VGND VPWR _1128_ _1131_ _1142_ _1130_ sg13g2_a21oi_1
XFILLER_7_394 VPWR VGND sg13g2_fill_2
X_4392_ _2083_ _2076_ _2079_ VPWR VGND sg13g2_nand2b_1
X_3343_ _1071_ VPWR _1073_ VGND _1041_ _1068_ sg13g2_o21ai_1
X_3274_ _1004_ net609 videogen.fancy_shader.n646\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_38_210 VPWR VGND sg13g2_decap_8
X_5013_ net118 VGND VPWR _0560_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\]
+ _0208_ sg13g2_dfrbpq_1
XFILLER_42_909 VPWR VGND sg13g2_decap_8
X_4962__371 VPWR VGND net371 sg13g2_tiehi
XFILLER_26_449 VPWR VGND sg13g2_decap_4
XFILLER_35_961 VPWR VGND sg13g2_fill_1
XFILLER_41_419 VPWR VGND sg13g2_decap_4
XFILLER_42_17 VPWR VGND sg13g2_fill_2
XFILLER_22_633 VPWR VGND sg13g2_decap_4
X_2989_ VGND VPWR _0832_ _0829_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ sg13g2_or2_1
X_4728_ net135 VGND VPWR _0279_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\]
+ _0010_ sg13g2_dfrbpq_1
X_4659_ net669 net719 _0212_ VPWR VGND sg13g2_nor2_1
XFILLER_18_917 VPWR VGND sg13g2_decap_8
XFILLER_29_243 VPWR VGND sg13g2_decap_8
XFILLER_44_202 VPWR VGND sg13g2_decap_4
XFILLER_16_51 VPWR VGND sg13g2_decap_4
XFILLER_26_961 VPWR VGND sg13g2_decap_8
XFILLER_41_942 VPWR VGND sg13g2_fill_1
XFILLER_41_986 VPWR VGND sg13g2_decap_8
XFILLER_12_121 VPWR VGND sg13g2_decap_8
XFILLER_13_666 VPWR VGND sg13g2_decap_8
XFILLER_12_165 VPWR VGND sg13g2_fill_1
XFILLER_12_176 VPWR VGND sg13g2_fill_1
X_4900__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_0_592 VPWR VGND sg13g2_fill_1
XFILLER_48_541 VPWR VGND sg13g2_decap_8
XFILLER_35_202 VPWR VGND sg13g2_fill_2
XFILLER_35_246 VPWR VGND sg13g2_decap_4
X_3961_ _1687_ net545 _1623_ VPWR VGND sg13g2_xnor2_1
X_2912_ _0703_ _0772_ _0787_ VPWR VGND sg13g2_nor2_2
X_3892_ _1619_ _1449_ _1616_ VPWR VGND sg13g2_nand2_1
XFILLER_31_441 VPWR VGND sg13g2_fill_2
X_2843_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\] net773 _0771_ _0418_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_997 VPWR VGND sg13g2_decap_8
X_2774_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\] _0755_ _0471_
+ VPWR VGND sg13g2_mux2_1
X_4513_ net675 net725 _0066_ VPWR VGND sg13g2_nor2_1
XFILLER_7_180 VPWR VGND sg13g2_fill_1
X_4444_ _2128_ VPWR _2133_ VGND _0646_ _2080_ sg13g2_o21ai_1
X_4375_ _2069_ tmds_green.dc_balancing_reg\[4\] _2068_ VPWR VGND sg13g2_xnor2_1
Xfanout605 tmds_blue.n100 net605 VPWR VGND sg13g2_buf_2
X_3326_ VPWR _1056_ net544 VGND sg13g2_inv_1
Xfanout627 net628 net627 VPWR VGND sg13g2_buf_8
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
Xfanout649 net650 net649 VPWR VGND sg13g2_buf_8
XFILLER_39_541 VPWR VGND sg13g2_decap_4
XFILLER_37_39 VPWR VGND sg13g2_fill_1
X_3257_ net747 _0992_ _0993_ _0364_ VPWR VGND sg13g2_nor3_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_3188_ _0949_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] _0948_ VPWR
+ VGND sg13g2_xnor2_1
XFILLER_23_920 VPWR VGND sg13g2_decap_8
XFILLER_23_997 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_fill_2
XFILLER_2_846 VPWR VGND sg13g2_decap_8
XFILLER_1_345 VPWR VGND sg13g2_decap_4
XFILLER_49_338 VPWR VGND sg13g2_decap_8
XFILLER_40_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_213 VPWR VGND sg13g2_fill_2
XFILLER_27_50 VPWR VGND sg13g2_fill_1
XFILLER_17_268 VPWR VGND sg13g2_fill_1
XFILLER_14_964 VPWR VGND sg13g2_decap_8
XFILLER_41_794 VPWR VGND sg13g2_fill_2
XFILLER_40_271 VPWR VGND sg13g2_decap_4
XFILLER_9_412 VPWR VGND sg13g2_fill_1
XFILLER_9_434 VPWR VGND sg13g2_fill_2
X_5022__35 VPWR VGND net35 sg13g2_tiehi
X_4802__370 VPWR VGND net370 sg13g2_tiehi
XFILLER_9_456 VPWR VGND sg13g2_fill_1
XFILLER_13_496 VPWR VGND sg13g2_fill_1
XFILLER_5_651 VPWR VGND sg13g2_fill_2
XFILLER_4_172 VPWR VGND sg13g2_decap_4
X_4160_ _1882_ VPWR _1883_ VGND _1876_ _1879_ sg13g2_o21ai_1
X_3111_ _0897_ _0791_ _0798_ _0896_ VPWR VGND sg13g2_and3_2
X_4091_ _1812_ _1731_ _1814_ VPWR VGND sg13g2_xor2_1
XFILLER_49_883 VPWR VGND sg13g2_decap_8
X_3042_ tmds_green.dc_balancing_reg\[0\] _0836_ _0263_ VPWR VGND sg13g2_and2_1
XFILLER_48_393 VPWR VGND sg13g2_decap_8
XFILLER_36_544 VPWR VGND sg13g2_decap_8
XFILLER_23_205 VPWR VGND sg13g2_decap_4
XFILLER_36_555 VPWR VGND sg13g2_fill_2
X_4993_ net223 VGND VPWR _0540_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\]
+ _0188_ sg13g2_dfrbpq_1
X_3944_ VGND VPWR _1662_ _1669_ _1670_ _1665_ sg13g2_a21oi_1
X_3875_ net623 _1600_ _1601_ _1603_ _1602_ net599 _1604_ VPWR VGND sg13g2_mux4_1
XFILLER_32_772 VPWR VGND sg13g2_decap_8
X_2826_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\] net753 _0768_ _0432_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_956 VPWR VGND sg13g2_decap_8
X_2757_ _0752_ _0715_ _0751_ VPWR VGND sg13g2_nand2_2
X_2688_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\] _0737_ _0548_
+ VPWR VGND sg13g2_mux2_1
X_4427_ _2106_ _2081_ _2109_ _2117_ VPWR VGND sg13g2_a21o_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_4358_ _2053_ tmds_green.dc_balancing_reg\[4\] _2052_ VPWR VGND sg13g2_xnor2_1
X_4289_ _1993_ _1989_ _1992_ VPWR VGND sg13g2_nand2_1
X_4884__228 VPWR VGND net228 sg13g2_tiehi
X_3309_ VPWR _1039_ _1038_ VGND sg13g2_inv_1
XFILLER_42_514 VPWR VGND sg13g2_fill_1
XFILLER_23_750 VPWR VGND sg13g2_decap_8
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_10_422 VPWR VGND sg13g2_decap_4
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_6_426 VPWR VGND sg13g2_fill_1
XFILLER_6_437 VPWR VGND sg13g2_fill_2
XFILLER_2_610 VPWR VGND sg13g2_decap_4
XFILLER_1_120 VPWR VGND sg13g2_fill_2
XFILLER_18_511 VPWR VGND sg13g2_fill_2
XFILLER_46_842 VPWR VGND sg13g2_decap_4
XFILLER_46_886 VPWR VGND sg13g2_decap_8
XFILLER_33_514 VPWR VGND sg13g2_fill_1
XFILLER_14_750 VPWR VGND sg13g2_decap_8
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_13_293 VPWR VGND sg13g2_fill_2
X_3660_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\] net561 _1390_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_253 VPWR VGND sg13g2_fill_1
XFILLER_9_264 VPWR VGND sg13g2_fill_2
X_2611_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\] _0711_ _0599_
+ VPWR VGND sg13g2_mux2_1
X_3591_ _1319_ _1320_ _1321_ VPWR VGND sg13g2_nor2_1
X_2542_ net413 net429 serialize.n433\[1\] VPWR VGND sg13g2_xor2_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_5_470 VPWR VGND sg13g2_fill_2
X_4212_ VGND VPWR _0642_ net607 _0497_ net750 sg13g2_a21oi_1
X_4143_ _1863_ _1862_ _1860_ _1866_ VPWR VGND sg13g2_a21o_1
X_4074_ _1010_ _1174_ _1797_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_319 VPWR VGND sg13g2_fill_1
X_3025_ net438 red_tmds_par\[0\] net698 serialize.n427\[0\] VPWR VGND sg13g2_mux2_1
XFILLER_11_208 VPWR VGND sg13g2_fill_1
X_4920__155 VPWR VGND net155 sg13g2_tiehi
X_4976_ net293 VGND VPWR _0523_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\]
+ _0171_ sg13g2_dfrbpq_1
X_3927_ _1635_ _1643_ _1647_ _1649_ _1653_ VPWR VGND sg13g2_nor4_1
XFILLER_20_720 VPWR VGND sg13g2_decap_8
Xclkload6 clknet_3_6__leaf_clk_regs clkload6/X VPWR VGND sg13g2_buf_1
X_3858_ net625 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\]
+ net628 _1587_ VPWR VGND sg13g2_mux4_1
XFILLER_30_1000 VPWR VGND sg13g2_decap_8
X_3789_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\] net550 _1519_ VPWR
+ VGND sg13g2_nor2_1
X_2809_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\] _0764_ _0445_
+ VPWR VGND sg13g2_mux2_1
XFILLER_4_908 VPWR VGND sg13g2_decap_8
XFILLER_46_149 VPWR VGND sg13g2_fill_1
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_28_886 VPWR VGND sg13g2_decap_8
XFILLER_27_363 VPWR VGND sg13g2_decap_8
XFILLER_11_720 VPWR VGND sg13g2_fill_2
XFILLER_7_702 VPWR VGND sg13g2_fill_2
XFILLER_10_230 VPWR VGND sg13g2_decap_4
XFILLER_10_252 VPWR VGND sg13g2_fill_2
XFILLER_40_83 VPWR VGND sg13g2_decap_4
XFILLER_3_974 VPWR VGND sg13g2_decap_8
XFILLER_2_440 VPWR VGND sg13g2_decap_4
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_37_138 VPWR VGND sg13g2_decap_8
XFILLER_1_66 VPWR VGND sg13g2_fill_1
XFILLER_46_694 VPWR VGND sg13g2_decap_4
XFILLER_19_886 VPWR VGND sg13g2_decap_4
X_4830_ net329 VGND VPWR _0381_ tmds_red.n114 net644 sg13g2_dfrbpq_2
XFILLER_21_528 VPWR VGND sg13g2_decap_4
X_4761_ net78 VGND VPWR _0312_ videogen.fancy_shader.video_x\[9\] net638 sg13g2_dfrbpq_2
XFILLER_14_1006 VPWR VGND sg13g2_decap_8
X_3712_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\] net556 _1442_ VPWR
+ VGND sg13g2_nor2_1
X_4692_ net684 net735 _0245_ VPWR VGND sg13g2_nor2_1
X_3643_ _1369_ _1370_ _1371_ _1372_ _1373_ VPWR VGND sg13g2_nor4_1
X_3574_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\] net555 _1304_ VPWR
+ VGND sg13g2_nor2_1
X_2525_ _0643_ net604 VPWR VGND sg13g2_inv_2
Xhold29 clockdiv.q0 VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold18 serialize.n411\[5\] VPWR VGND net423 sg13g2_dlygate4sd3_1
X_4126_ _1837_ _1847_ _1831_ _1849_ VPWR VGND sg13g2_nand3_1
XFILLER_29_617 VPWR VGND sg13g2_decap_8
X_4057_ _1780_ _1778_ _1779_ VPWR VGND sg13g2_nand2b_1
X_3008_ net443 blue_tmds_par\[2\] net695 serialize.n429\[4\] VPWR VGND sg13g2_mux2_1
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_25_823 VPWR VGND sg13g2_decap_8
XFILLER_25_878 VPWR VGND sg13g2_decap_8
XFILLER_24_366 VPWR VGND sg13g2_decap_4
X_4959_ net383 VGND VPWR _0506_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\]
+ _0154_ sg13g2_dfrbpq_1
XFILLER_0_933 VPWR VGND sg13g2_decap_8
XFILLER_48_937 VPWR VGND sg13g2_decap_8
XFILLER_47_425 VPWR VGND sg13g2_decap_8
XFILLER_16_823 VPWR VGND sg13g2_decap_8
XFILLER_27_160 VPWR VGND sg13g2_fill_2
XFILLER_27_171 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_fill_1
XFILLER_42_163 VPWR VGND sg13g2_fill_1
XFILLER_31_804 VPWR VGND sg13g2_decap_8
XFILLER_35_72 VPWR VGND sg13g2_fill_1
XFILLER_31_837 VPWR VGND sg13g2_decap_8
XFILLER_30_358 VPWR VGND sg13g2_decap_4
XFILLER_7_587 VPWR VGND sg13g2_fill_2
X_3290_ VGND VPWR _1020_ _1018_ _1010_ sg13g2_or2_1
XFILLER_39_937 VPWR VGND sg13g2_fill_1
XFILLER_39_926 VPWR VGND sg13g2_decap_8
X_4910__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_19_650 VPWR VGND sg13g2_decap_4
XFILLER_34_653 VPWR VGND sg13g2_fill_1
X_4813_ net348 VGND VPWR _0364_ videogen.fancy_shader.video_y\[8\] net635 sg13g2_dfrbpq_2
X_4744_ net103 VGND VPWR _0295_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\]
+ _0026_ sg13g2_dfrbpq_1
XFILLER_30_881 VPWR VGND sg13g2_decap_8
XFILLER_31_19 VPWR VGND sg13g2_fill_2
X_4675_ net686 net737 _0228_ VPWR VGND sg13g2_nor2_1
X_3626_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\] net565 _1356_ VPWR
+ VGND sg13g2_nor2_1
Xoutput19 net19 uo_out[6] VPWR VGND sg13g2_buf_1
X_3557_ net597 _1281_ _1286_ _1287_ VPWR VGND sg13g2_nor3_1
X_3488_ _1037_ _1211_ _1218_ VPWR VGND sg13g2_and2_1
XFILLER_45_929 VPWR VGND sg13g2_decap_8
X_5089_ net798 VGND VPWR serialize.n428\[4\] serialize.n414\[2\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4109_ _1803_ _1826_ _1830_ _1832_ VPWR VGND sg13g2_or3_1
XFILLER_25_642 VPWR VGND sg13g2_decap_8
XFILLER_25_686 VPWR VGND sg13g2_decap_8
XFILLER_21_870 VPWR VGND sg13g2_decap_8
XFILLER_4_579 VPWR VGND sg13g2_decap_4
XFILLER_0_730 VPWR VGND sg13g2_decap_8
XFILLER_46_60 VPWR VGND sg13g2_decap_4
XFILLER_29_981 VPWR VGND sg13g2_decap_8
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_43_461 VPWR VGND sg13g2_decap_8
XFILLER_7_10 VPWR VGND sg13g2_fill_2
X_2790_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\] net778 _0758_ _0458_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_852 VPWR VGND sg13g2_fill_2
X_4460_ net651 net702 _0013_ VPWR VGND sg13g2_nor2_1
X_4391_ _2082_ tmds_blue.dc_balancing_reg\[2\] _2080_ VPWR VGND sg13g2_xnor2_1
X_3411_ _1138_ _1139_ _1136_ _1141_ VPWR VGND sg13g2_nand3_1
X_3342_ _1072_ _1070_ _1057_ _1069_ _1042_ VPWR VGND sg13g2_a22oi_1
X_4812__350 VPWR VGND net350 sg13g2_tiehi
X_3273_ _1003_ net608 videogen.fancy_shader.n646\[1\] VPWR VGND sg13g2_nand2_1
X_5012_ net126 VGND VPWR _0559_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\]
+ _0207_ sg13g2_dfrbpq_1
XFILLER_35_984 VPWR VGND sg13g2_decap_8
XFILLER_22_645 VPWR VGND sg13g2_decap_8
X_2988_ _0820_ _0831_ net20 VPWR VGND sg13g2_nor2_1
X_4727_ net136 VGND VPWR _0278_ red_tmds_par\[7\] net645 sg13g2_dfrbpq_1
X_4658_ net684 net719 _0211_ VPWR VGND sg13g2_nor2_1
X_3609_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\] net575 _1339_ VPWR
+ VGND sg13g2_nor2_1
X_4589_ net687 net738 _0142_ VPWR VGND sg13g2_nor2_1
XFILLER_44_214 VPWR VGND sg13g2_fill_1
XFILLER_29_266 VPWR VGND sg13g2_decap_8
XFILLER_45_759 VPWR VGND sg13g2_fill_1
XFILLER_26_940 VPWR VGND sg13g2_decap_8
XFILLER_41_965 VPWR VGND sg13g2_decap_8
X_4894__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_9_616 VPWR VGND sg13g2_decap_8
XFILLER_13_656 VPWR VGND sg13g2_fill_2
XFILLER_8_126 VPWR VGND sg13g2_fill_1
XFILLER_32_40 VPWR VGND sg13g2_fill_1
XFILLER_12_188 VPWR VGND sg13g2_decap_4
XFILLER_32_84 VPWR VGND sg13g2_fill_1
XFILLER_32_95 VPWR VGND sg13g2_fill_2
X_4794__386 VPWR VGND net386 sg13g2_tiehi
XFILLER_48_520 VPWR VGND sg13g2_decap_8
XFILLER_48_597 VPWR VGND sg13g2_decap_8
XFILLER_17_984 VPWR VGND sg13g2_decap_8
X_3960_ _1684_ _1685_ _1686_ VPWR VGND sg13g2_and2_1
XFILLER_44_792 VPWR VGND sg13g2_fill_1
XFILLER_16_494 VPWR VGND sg13g2_fill_1
X_2911_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\] _0786_ _0291_
+ VPWR VGND sg13g2_mux2_1
XFILLER_43_291 VPWR VGND sg13g2_decap_4
X_3891_ VGND VPWR _1351_ _1618_ _0373_ _1551_ sg13g2_a21oi_1
XFILLER_32_976 VPWR VGND sg13g2_decap_8
X_2842_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\] net768 _0771_ _0419_
+ VPWR VGND sg13g2_mux2_1
X_2773_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\] _0755_ _0472_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_671 VPWR VGND sg13g2_fill_2
X_4512_ net674 net726 _0065_ VPWR VGND sg13g2_nor2_1
XFILLER_7_170 VPWR VGND sg13g2_decap_4
X_4443_ _2131_ VPWR _2132_ VGND _2097_ _2119_ sg13g2_o21ai_1
X_4374_ _2024_ VPWR _2068_ VGND _0641_ _2022_ sg13g2_o21ai_1
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
Xfanout628 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[0\] net628 VPWR VGND
+ sg13g2_buf_8
X_3325_ _1055_ _1053_ _1054_ VPWR VGND sg13g2_nand2_2
Xfanout639 net650 net639 VPWR VGND sg13g2_buf_2
Xfanout617 net618 net617 VPWR VGND sg13g2_buf_2
X_3256_ videogen.fancy_shader.video_y\[8\] _0991_ _0993_ VPWR VGND sg13g2_and2_1
XFILLER_39_575 VPWR VGND sg13g2_decap_8
XFILLER_2_1007 VPWR VGND sg13g2_decap_8
X_3187_ _0915_ _0919_ _0947_ _0948_ _0331_ VPWR VGND sg13g2_nor4_1
XFILLER_27_715 VPWR VGND sg13g2_decap_8
XFILLER_26_236 VPWR VGND sg13g2_decap_8
XFILLER_35_770 VPWR VGND sg13g2_fill_2
XFILLER_23_976 VPWR VGND sg13g2_decap_8
XFILLER_6_619 VPWR VGND sg13g2_decap_8
XFILLER_5_129 VPWR VGND sg13g2_decap_4
XFILLER_2_825 VPWR VGND sg13g2_decap_8
XFILLER_49_317 VPWR VGND sg13g2_decap_8
XFILLER_18_759 VPWR VGND sg13g2_decap_8
XFILLER_26_792 VPWR VGND sg13g2_fill_1
XFILLER_13_420 VPWR VGND sg13g2_fill_1
XFILLER_14_943 VPWR VGND sg13g2_decap_8
XFILLER_25_280 VPWR VGND sg13g2_decap_8
XFILLER_43_61 VPWR VGND sg13g2_decap_8
XFILLER_5_685 VPWR VGND sg13g2_fill_1
XFILLER_4_195 VPWR VGND sg13g2_decap_8
X_3110_ net629 videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\]
+ _0896_ VPWR VGND sg13g2_nor3_1
X_4090_ _1813_ _1731_ _1812_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_390 VPWR VGND sg13g2_fill_2
XFILLER_49_862 VPWR VGND sg13g2_decap_8
X_3041_ _0837_ net606 net796 VPWR VGND sg13g2_nand2_1
XFILLER_48_372 VPWR VGND sg13g2_decap_8
XFILLER_36_578 VPWR VGND sg13g2_fill_1
X_4992_ net227 VGND VPWR _0539_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\]
+ _0187_ sg13g2_dfrbpq_1
X_3943_ _1667_ _1668_ _1669_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_935 VPWR VGND sg13g2_decap_8
X_3874_ net624 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\]
+ net627 _1603_ VPWR VGND sg13g2_mux4_1
X_2825_ _0723_ _0762_ _0768_ VPWR VGND sg13g2_nor2_2
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_2756_ _0679_ _0705_ _0751_ VPWR VGND sg13g2_nor2_2
X_2687_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\] _0737_ _0549_
+ VPWR VGND sg13g2_mux2_1
X_4426_ _2106_ _2109_ _2081_ _2116_ VPWR VGND sg13g2_nand3_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4357_ VGND VPWR tmds_green.dc_balancing_reg\[3\] _2024_ _2052_ _2022_ sg13g2_a21oi_1
X_4288_ _1992_ _0643_ _1991_ VPWR VGND sg13g2_xnor2_1
X_3308_ _1016_ _1025_ _1038_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_309 VPWR VGND sg13g2_decap_8
X_3239_ _0982_ videogen.fancy_shader.video_y\[2\] _0976_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_504 VPWR VGND sg13g2_decap_4
XFILLER_42_537 VPWR VGND sg13g2_fill_1
XFILLER_42_526 VPWR VGND sg13g2_decap_8
XFILLER_23_784 VPWR VGND sg13g2_decap_8
XFILLER_11_935 VPWR VGND sg13g2_decap_8
XFILLER_6_416 VPWR VGND sg13g2_fill_2
XFILLER_6_449 VPWR VGND sg13g2_decap_4
XFILLER_2_622 VPWR VGND sg13g2_fill_2
XFILLER_1_187 VPWR VGND sg13g2_decap_8
XFILLER_46_810 VPWR VGND sg13g2_decap_8
XFILLER_37_309 VPWR VGND sg13g2_decap_4
XFILLER_46_832 VPWR VGND sg13g2_fill_1
XFILLER_46_821 VPWR VGND sg13g2_fill_2
XFILLER_46_865 VPWR VGND sg13g2_decap_8
XFILLER_45_397 VPWR VGND sg13g2_fill_1
XFILLER_33_526 VPWR VGND sg13g2_decap_8
XFILLER_9_276 VPWR VGND sg13g2_decap_8
X_3590_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\] net561 _1320_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_287 VPWR VGND sg13g2_decap_8
X_2610_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\] _0711_ _0600_
+ VPWR VGND sg13g2_mux2_1
X_2541_ _0658_ net429 net413 VPWR VGND sg13g2_nand2_1
XFILLER_5_482 VPWR VGND sg13g2_fill_2
X_4211_ net751 _1924_ _0388_ VPWR VGND sg13g2_nor2_1
X_4142_ VGND VPWR _1862_ _1863_ _1865_ _1860_ sg13g2_a21oi_1
XFILLER_37_810 VPWR VGND sg13g2_fill_2
X_4073_ _1725_ _1174_ _1796_ VPWR VGND sg13g2_xor2_1
X_3024_ green_tmds_par\[9\] net699 serialize.n428\[9\] VPWR VGND sg13g2_and2_1
XFILLER_37_832 VPWR VGND sg13g2_fill_2
XFILLER_37_821 VPWR VGND sg13g2_decap_8
XFILLER_37_876 VPWR VGND sg13g2_fill_2
XFILLER_24_515 VPWR VGND sg13g2_fill_1
X_4975_ net297 VGND VPWR _0522_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\]
+ _0170_ sg13g2_dfrbpq_1
X_3926_ _1652_ _1634_ _1650_ VPWR VGND sg13g2_nand2_1
Xclkload7 VPWR clkload7/Y clknet_3_7__leaf_clk_regs VGND sg13g2_inv_1
X_3857_ net620 VPWR _1586_ VGND _1568_ _1585_ sg13g2_o21ai_1
X_3788_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\] net560 _1518_ VPWR
+ VGND sg13g2_nor2_1
X_2808_ net778 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\] _0764_ _0446_
+ VPWR VGND sg13g2_mux2_1
X_2739_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\] _0747_ _0507_
+ VPWR VGND sg13g2_mux2_1
X_4409_ VGND VPWR net604 _2074_ _2100_ _2088_ sg13g2_a21oi_1
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
XFILLER_47_618 VPWR VGND sg13g2_decap_8
X_5027__349 VPWR VGND net349 sg13g2_tiehi
XFILLER_28_854 VPWR VGND sg13g2_fill_1
XFILLER_15_548 VPWR VGND sg13g2_fill_1
XFILLER_3_953 VPWR VGND sg13g2_decap_8
XFILLER_34_9 VPWR VGND sg13g2_decap_4
XFILLER_33_301 VPWR VGND sg13g2_fill_1
X_5004__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_33_334 VPWR VGND sg13g2_decap_8
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_34_879 VPWR VGND sg13g2_decap_8
X_4760_ net79 VGND VPWR _0311_ videogen.fancy_shader.video_x\[8\] net638 sg13g2_dfrbpq_2
X_3711_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\] net589 _1441_ VPWR
+ VGND sg13g2_nor2_1
X_4691_ net684 net735 _0244_ VPWR VGND sg13g2_nor2_1
X_3642_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\] net575 _1372_ VPWR
+ VGND sg13g2_nor2_1
X_3573_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\] net565 _1303_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2524_ _0642_ tmds_green.dc_balancing_reg\[4\] VPWR VGND sg13g2_inv_2
XFILLER_29_19 VPWR VGND sg13g2_fill_2
Xhold19 serialize.n411\[7\] VPWR VGND net424 sg13g2_dlygate4sd3_1
X_4125_ _1837_ _1831_ _1847_ _1848_ VPWR VGND sg13g2_a21o_1
XFILLER_28_139 VPWR VGND sg13g2_fill_2
X_4056_ _1779_ _1688_ _1725_ VPWR VGND sg13g2_xnor2_1
X_3007_ net436 blue_tmds_par\[3\] net695 serialize.n429\[3\] VPWR VGND sg13g2_mux2_1
XFILLER_36_183 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_4
X_4958_ net385 VGND VPWR _0505_ tmds_red.dc_balancing_reg\[4\] net647 sg13g2_dfrbpq_2
X_4889_ net218 VGND VPWR _0440_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\]
+ _0097_ sg13g2_dfrbpq_1
X_3909_ _1635_ _1634_ VPWR VGND sg13g2_inv_2
XFILLER_20_573 VPWR VGND sg13g2_decap_8
XFILLER_3_238 VPWR VGND sg13g2_fill_2
XFILLER_0_912 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_fill_1
XFILLER_48_916 VPWR VGND sg13g2_decap_8
XFILLER_0_989 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_fill_1
XFILLER_15_312 VPWR VGND sg13g2_fill_1
XFILLER_37_1018 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_24_890 VPWR VGND sg13g2_decap_8
X_5073__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_11_540 VPWR VGND sg13g2_fill_1
XFILLER_11_551 VPWR VGND sg13g2_decap_8
XFILLER_7_533 VPWR VGND sg13g2_fill_2
XFILLER_7_555 VPWR VGND sg13g2_decap_8
X_5010__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_2_293 VPWR VGND sg13g2_fill_2
XFILLER_38_415 VPWR VGND sg13g2_fill_2
XFILLER_18_183 VPWR VGND sg13g2_fill_1
X_4812_ net350 VGND VPWR _0363_ videogen.fancy_shader.video_y\[7\] net636 sg13g2_dfrbpq_2
XFILLER_22_838 VPWR VGND sg13g2_decap_8
XFILLER_33_197 VPWR VGND sg13g2_decap_8
X_4743_ net105 VGND VPWR _0294_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\]
+ _0025_ sg13g2_dfrbpq_1
X_4674_ net671 net723 _0227_ VPWR VGND sg13g2_nor2_1
X_3625_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\] net588 _1355_ VPWR
+ VGND sg13g2_nor2_1
X_3556_ _1282_ _1283_ _1284_ _1285_ _1286_ VPWR VGND sg13g2_nor4_1
X_4735__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_0_219 VPWR VGND sg13g2_decap_8
X_3487_ VGND VPWR _1211_ _1216_ _1217_ _1037_ sg13g2_a21oi_1
XFILLER_5_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_1016 VPWR VGND sg13g2_decap_8
XFILLER_45_908 VPWR VGND sg13g2_decap_8
X_5088_ net801 VGND VPWR serialize.n428\[3\] serialize.n414\[1\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4108_ _1803_ _1830_ _1831_ VPWR VGND sg13g2_nor2_1
XFILLER_29_459 VPWR VGND sg13g2_decap_4
XFILLER_44_407 VPWR VGND sg13g2_fill_1
XFILLER_38_993 VPWR VGND sg13g2_decap_8
X_4039_ VPWR VGND _1752_ _1757_ _1756_ _1749_ _1762_ _1753_ sg13g2_a221oi_1
XFILLER_24_164 VPWR VGND sg13g2_decap_8
XFILLER_12_337 VPWR VGND sg13g2_fill_2
XFILLER_0_786 VPWR VGND sg13g2_decap_8
XFILLER_29_960 VPWR VGND sg13g2_decap_8
XFILLER_35_407 VPWR VGND sg13g2_fill_2
XFILLER_28_481 VPWR VGND sg13g2_decap_8
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_15_142 VPWR VGND sg13g2_decap_4
XFILLER_15_153 VPWR VGND sg13g2_decap_8
XFILLER_31_668 VPWR VGND sg13g2_decap_8
XFILLER_8_831 VPWR VGND sg13g2_fill_1
XFILLER_8_820 VPWR VGND sg13g2_decap_8
X_4945__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_30_167 VPWR VGND sg13g2_decap_8
X_4955__391 VPWR VGND net391 sg13g2_tiehi
X_4390_ _2081_ _2080_ tmds_blue.dc_balancing_reg\[2\] VPWR VGND sg13g2_nand2b_1
X_3410_ _1138_ _1139_ _1140_ VPWR VGND sg13g2_and2_1
X_3341_ _1071_ _1057_ _1070_ VPWR VGND sg13g2_nand2_1
X_3272_ net748 _1002_ _0370_ VPWR VGND sg13g2_nor2_1
X_5011_ net134 VGND VPWR _0558_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\]
+ _0206_ sg13g2_dfrbpq_1
XFILLER_27_919 VPWR VGND sg13g2_decap_8
XFILLER_35_930 VPWR VGND sg13g2_fill_1
XFILLER_42_19 VPWR VGND sg13g2_fill_1
X_2987_ VGND VPWR _0829_ _0830_ _0831_ _0819_ sg13g2_a21oi_1
X_4726_ net137 VGND VPWR _0277_ red_tmds_par\[5\] net645 sg13g2_dfrbpq_1
X_4657_ net669 net719 _0210_ VPWR VGND sg13g2_nor2_1
X_3608_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\] net551 _1338_ VPWR
+ VGND sg13g2_nor2_1
X_4588_ net677 net729 _0141_ VPWR VGND sg13g2_nor2_1
X_3539_ _1265_ _1266_ _1267_ _1268_ _1269_ VPWR VGND sg13g2_nor4_1
XFILLER_27_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_223 VPWR VGND sg13g2_fill_1
XFILLER_44_259 VPWR VGND sg13g2_fill_2
XFILLER_25_451 VPWR VGND sg13g2_fill_2
XFILLER_41_933 VPWR VGND sg13g2_decap_8
XFILLER_13_602 VPWR VGND sg13g2_fill_2
XFILLER_25_484 VPWR VGND sg13g2_fill_2
XFILLER_26_996 VPWR VGND sg13g2_decap_8
XFILLER_40_487 VPWR VGND sg13g2_fill_2
XFILLER_8_138 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_fill_2
X_5070__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_4_333 VPWR VGND sg13g2_decap_4
XFILLER_4_311 VPWR VGND sg13g2_fill_1
XFILLER_10_1010 VPWR VGND sg13g2_decap_8
XFILLER_0_583 VPWR VGND sg13g2_decap_8
XFILLER_48_576 VPWR VGND sg13g2_decap_8
X_5042__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_36_705 VPWR VGND sg13g2_fill_2
XFILLER_17_963 VPWR VGND sg13g2_decap_8
XFILLER_43_270 VPWR VGND sg13g2_decap_8
X_2910_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\] _0786_ _0292_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_484 VPWR VGND sg13g2_fill_2
X_3890_ _1551_ _1618_ _0374_ VPWR VGND sg13g2_nor2_1
XFILLER_31_443 VPWR VGND sg13g2_fill_1
XFILLER_32_955 VPWR VGND sg13g2_decap_8
X_2841_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\] net753 _0771_ _0420_
+ VPWR VGND sg13g2_mux2_1
X_2772_ _0755_ _0717_ _0751_ VPWR VGND sg13g2_nand2_2
XFILLER_8_650 VPWR VGND sg13g2_decap_8
X_4511_ net675 net725 _0064_ VPWR VGND sg13g2_nor2_1
X_4442_ _2131_ _2127_ _2130_ VPWR VGND sg13g2_xnor2_1
X_4373_ _2057_ _2066_ _2067_ VPWR VGND sg13g2_nor2_1
Xfanout629 videogen.fancy_shader.video_x\[7\] net629 VPWR VGND sg13g2_buf_8
X_3324_ _1054_ _1046_ _1052_ VPWR VGND sg13g2_nand2_1
Xfanout607 display_enable net607 VPWR VGND sg13g2_buf_8
Xfanout618 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net618 VPWR VGND
+ sg13g2_buf_8
X_3255_ videogen.fancy_shader.video_y\[8\] _0991_ _0992_ VPWR VGND sg13g2_nor2_1
X_3186_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\] _0946_ _0948_ VPWR
+ VGND sg13g2_and2_1
X_4923__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_41_229 VPWR VGND sg13g2_decap_8
XFILLER_22_421 VPWR VGND sg13g2_fill_2
XFILLER_23_955 VPWR VGND sg13g2_decap_8
XFILLER_34_292 VPWR VGND sg13g2_fill_1
XFILLER_10_616 VPWR VGND sg13g2_decap_8
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_108 VPWR VGND sg13g2_fill_2
X_4709_ net656 net707 _0260_ VPWR VGND sg13g2_nor2_1
X_4932__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_45_535 VPWR VGND sg13g2_decap_8
XFILLER_17_215 VPWR VGND sg13g2_fill_1
XFILLER_14_922 VPWR VGND sg13g2_decap_8
XFILLER_26_760 VPWR VGND sg13g2_fill_2
XFILLER_13_443 VPWR VGND sg13g2_fill_1
XFILLER_13_476 VPWR VGND sg13g2_decap_8
XFILLER_14_999 VPWR VGND sg13g2_decap_8
XFILLER_9_436 VPWR VGND sg13g2_fill_1
XFILLER_5_653 VPWR VGND sg13g2_fill_1
XFILLER_1_881 VPWR VGND sg13g2_decap_8
XFILLER_49_841 VPWR VGND sg13g2_decap_8
XFILLER_48_351 VPWR VGND sg13g2_decap_8
X_3040_ _0647_ net750 _0836_ VPWR VGND sg13g2_nor2_2
XFILLER_24_719 VPWR VGND sg13g2_decap_8
X_4991_ net231 VGND VPWR _0538_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\]
+ _0186_ sg13g2_dfrbpq_1
X_3942_ _1645_ _1654_ _1668_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_914 VPWR VGND sg13g2_decap_8
X_3873_ net627 videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\]
+ net624 _1602_ VPWR VGND sg13g2_mux4_1
X_2824_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\] net788 _0767_ _0433_
+ VPWR VGND sg13g2_mux2_1
X_2755_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\] _0750_ _0485_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_480 VPWR VGND sg13g2_fill_1
X_4772__58 VPWR VGND net58 sg13g2_tiehi
X_2686_ _0737_ _0717_ _0720_ VPWR VGND sg13g2_nand2_2
X_4425_ VPWR _2115_ _2114_ VGND sg13g2_inv_1
X_4356_ VGND VPWR _2046_ _2048_ _2051_ _2045_ sg13g2_a21oi_1
X_4853__292 VPWR VGND net292 sg13g2_tiehi
X_3307_ VPWR _1037_ _1036_ VGND sg13g2_inv_1
XFILLER_24_1009 VPWR VGND sg13g2_decap_8
X_4287_ _1990_ VPWR _1991_ VGND tmds_blue.n193 _0644_ sg13g2_o21ai_1
XFILLER_39_340 VPWR VGND sg13g2_fill_2
X_3238_ _0981_ net795 _0980_ VPWR VGND sg13g2_nand2_1
X_3169_ _0793_ _0935_ _0936_ _0325_ VPWR VGND sg13g2_nor3_1
XFILLER_15_708 VPWR VGND sg13g2_decap_8
XFILLER_15_719 VPWR VGND sg13g2_fill_1
XFILLER_27_546 VPWR VGND sg13g2_fill_2
XFILLER_27_579 VPWR VGND sg13g2_decap_8
XFILLER_35_590 VPWR VGND sg13g2_fill_1
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_13_43 VPWR VGND sg13g2_fill_2
XFILLER_1_122 VPWR VGND sg13g2_fill_1
X_4715__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_49_148 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_4
XFILLER_18_513 VPWR VGND sg13g2_fill_1
XFILLER_46_855 VPWR VGND sg13g2_fill_1
X_2540_ VPWR _0657_ net421 VGND sg13g2_inv_1
XFILLER_6_984 VPWR VGND sg13g2_decap_8
X_4210_ _0647_ _0891_ _1924_ VPWR VGND sg13g2_nor2_1
X_4141_ _1864_ _1862_ _1863_ VPWR VGND sg13g2_nand2_1
X_4072_ _1792_ _1794_ _1791_ _1795_ VPWR VGND sg13g2_nand3_1
X_3023_ green_tmds_par\[8\] net696 serialize.n428\[8\] VPWR VGND sg13g2_and2_1
X_4883__230 VPWR VGND net230 sg13g2_tiehi
X_4809__356 VPWR VGND net356 sg13g2_tiehi
XFILLER_36_332 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
X_4974_ net300 VGND VPWR _0521_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\]
+ _0169_ sg13g2_dfrbpq_1
XFILLER_17_590 VPWR VGND sg13g2_decap_8
X_3925_ VPWR _1651_ _1650_ VGND sg13g2_inv_1
X_3856_ _1566_ VPWR _1585_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\]
+ net550 sg13g2_o21ai_1
X_3787_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\] net573 _1517_ VPWR
+ VGND sg13g2_nor2_1
X_2807_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\] _0764_ _0447_
+ VPWR VGND sg13g2_mux2_1
X_2738_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\] _0747_ _0508_
+ VPWR VGND sg13g2_mux2_1
X_4408_ _2002_ _2098_ _2099_ VPWR VGND sg13g2_nor2_1
X_2669_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\] _0733_ _0563_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
X_4786__404 VPWR VGND net404 sg13g2_tiehi
X_4339_ _2035_ _2033_ _2029_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_170 VPWR VGND sg13g2_fill_1
XFILLER_39_181 VPWR VGND sg13g2_decap_4
X_4745__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_42_324 VPWR VGND sg13g2_decap_8
XFILLER_11_744 VPWR VGND sg13g2_fill_1
XFILLER_7_759 VPWR VGND sg13g2_decap_4
XFILLER_10_254 VPWR VGND sg13g2_fill_1
XFILLER_10_265 VPWR VGND sg13g2_fill_1
XFILLER_11_799 VPWR VGND sg13g2_decap_4
XFILLER_40_30 VPWR VGND sg13g2_fill_1
XFILLER_6_236 VPWR VGND sg13g2_fill_1
XFILLER_10_287 VPWR VGND sg13g2_decap_8
XFILLER_3_932 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_decap_8
XFILLER_38_608 VPWR VGND sg13g2_decap_8
XFILLER_37_118 VPWR VGND sg13g2_fill_2
XFILLER_19_822 VPWR VGND sg13g2_fill_2
Xfanout790 net791 net790 VPWR VGND sg13g2_buf_8
XFILLER_33_313 VPWR VGND sg13g2_decap_8
XFILLER_34_858 VPWR VGND sg13g2_decap_8
XFILLER_42_891 VPWR VGND sg13g2_decap_8
XFILLER_14_571 VPWR VGND sg13g2_decap_8
XFILLER_14_593 VPWR VGND sg13g2_decap_8
X_3710_ net597 VPWR _1440_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\]
+ net567 sg13g2_o21ai_1
X_4690_ net685 net736 _0243_ VPWR VGND sg13g2_nor2_1
X_3641_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\] net551 _1371_ VPWR
+ VGND sg13g2_nor2_1
X_3572_ net622 VPWR _1302_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\]
+ net588 sg13g2_o21ai_1
X_2523_ VPWR _0641_ tmds_green.dc_balancing_reg\[3\] VGND sg13g2_inv_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_4124_ _1833_ _1846_ _1847_ VPWR VGND sg13g2_nor2b_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_2
XFILLER_28_107 VPWR VGND sg13g2_fill_2
XFILLER_49_490 VPWR VGND sg13g2_decap_8
X_4055_ _1776_ _1773_ _1778_ VPWR VGND sg13g2_xor2_1
X_3006_ net441 blue_tmds_par\[2\] net695 serialize.n429\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_37_674 VPWR VGND sg13g2_decap_8
XFILLER_25_836 VPWR VGND sg13g2_decap_4
XFILLER_25_847 VPWR VGND sg13g2_fill_2
XFILLER_40_828 VPWR VGND sg13g2_fill_2
XFILLER_40_817 VPWR VGND sg13g2_decap_8
XFILLER_24_379 VPWR VGND sg13g2_decap_8
X_4957_ net387 VGND VPWR _0504_ tmds_red.dc_balancing_reg\[3\] net647 sg13g2_dfrbpq_1
XFILLER_33_891 VPWR VGND sg13g2_decap_4
X_3908_ _1633_ _1060_ _1634_ VPWR VGND sg13g2_xor2_1
X_4888_ net220 VGND VPWR _0439_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\]
+ _0096_ sg13g2_dfrbpq_1
X_3839_ _1567_ VPWR _1568_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\]
+ net560 sg13g2_o21ai_1
XFILLER_4_729 VPWR VGND sg13g2_decap_8
XFILLER_0_968 VPWR VGND sg13g2_decap_8
XFILLER_16_836 VPWR VGND sg13g2_decap_8
XFILLER_43_666 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_fill_2
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_43_699 VPWR VGND sg13g2_decap_4
XFILLER_42_187 VPWR VGND sg13g2_decap_8
XFILLER_30_316 VPWR VGND sg13g2_fill_1
XFILLER_42_198 VPWR VGND sg13g2_fill_2
XFILLER_3_740 VPWR VGND sg13g2_fill_1
XFILLER_2_272 VPWR VGND sg13g2_decap_8
XFILLER_2_283 VPWR VGND sg13g2_fill_2
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_46_493 VPWR VGND sg13g2_fill_2
XFILLER_34_644 VPWR VGND sg13g2_decap_8
X_4811_ net352 VGND VPWR _0362_ videogen.fancy_shader.video_y\[6\] net635 sg13g2_dfrbpq_2
XFILLER_22_817 VPWR VGND sg13g2_decap_8
XFILLER_33_176 VPWR VGND sg13g2_fill_2
X_4742_ net107 VGND VPWR _0293_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\]
+ _0024_ sg13g2_dfrbpq_1
X_4673_ net686 net738 _0226_ VPWR VGND sg13g2_nor2_1
X_3624_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\] net555 _1354_ VPWR
+ VGND sg13g2_nor2_1
X_3555_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\] net587 _1285_ VPWR
+ VGND sg13g2_nor2_1
X_3486_ _1204_ _1212_ _1036_ _1216_ VPWR VGND _1214_ sg13g2_nand4_1
XFILLER_29_416 VPWR VGND sg13g2_fill_2
X_5087_ net799 VGND VPWR serialize.n428\[2\] serialize.n414\[0\] clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_38_950 VPWR VGND sg13g2_decap_8
X_4107_ _1830_ _1806_ _1829_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_972 VPWR VGND sg13g2_decap_8
X_4038_ _1761_ _1758_ _1760_ _1753_ _1749_ VPWR VGND sg13g2_a22oi_1
XFILLER_40_658 VPWR VGND sg13g2_decap_4
XFILLER_12_349 VPWR VGND sg13g2_decap_8
XFILLER_20_360 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_4
XFILLER_43_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_765 VPWR VGND sg13g2_decap_8
XFILLER_48_747 VPWR VGND sg13g2_decap_8
XFILLER_28_460 VPWR VGND sg13g2_fill_1
XFILLER_46_95 VPWR VGND sg13g2_decap_4
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_43_430 VPWR VGND sg13g2_decap_4
XFILLER_16_666 VPWR VGND sg13g2_decap_8
XFILLER_31_614 VPWR VGND sg13g2_decap_8
XFILLER_7_12 VPWR VGND sg13g2_fill_1
XFILLER_7_331 VPWR VGND sg13g2_decap_4
XFILLER_11_382 VPWR VGND sg13g2_decap_4
XFILLER_8_898 VPWR VGND sg13g2_decap_8
X_3340_ _1043_ VPWR _1070_ VGND _0634_ _0640_ sg13g2_o21ai_1
XFILLER_3_581 VPWR VGND sg13g2_decap_8
X_3271_ VGND VPWR _0668_ _0797_ _1002_ _1001_ sg13g2_a21oi_1
X_5010_ net150 VGND VPWR _0557_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\]
+ _0205_ sg13g2_dfrbpq_1
XFILLER_39_769 VPWR VGND sg13g2_fill_2
XFILLER_38_235 VPWR VGND sg13g2_fill_2
XFILLER_38_224 VPWR VGND sg13g2_decap_8
XFILLER_19_471 VPWR VGND sg13g2_fill_2
X_2986_ _0825_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\]
+ _0830_ VPWR VGND sg13g2_a21o_1
X_4725_ net138 VGND VPWR _0276_ red_tmds_par\[3\] net645 sg13g2_dfrbpq_1
X_4656_ net669 net719 _0209_ VPWR VGND sg13g2_nor2_1
X_5030__302 VPWR VGND net302 sg13g2_tiehi
X_4587_ net676 net729 _0140_ VPWR VGND sg13g2_nor2_1
X_3607_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\] net585 _1337_ VPWR
+ VGND sg13g2_nor2_1
X_3538_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\] net553 _1268_ VPWR
+ VGND sg13g2_nor2_1
X_3469_ VPWR VGND _1191_ _1196_ _1190_ _1085_ _1199_ _1086_ sg13g2_a221oi_1
XFILLER_44_238 VPWR VGND sg13g2_fill_1
X_4863__272 VPWR VGND net272 sg13g2_tiehi
XFILLER_26_975 VPWR VGND sg13g2_decap_8
XFILLER_16_87 VPWR VGND sg13g2_fill_1
XFILLER_13_658 VPWR VGND sg13g2_fill_1
XFILLER_21_691 VPWR VGND sg13g2_fill_2
XFILLER_5_813 VPWR VGND sg13g2_decap_4
XFILLER_32_97 VPWR VGND sg13g2_fill_1
XFILLER_48_500 VPWR VGND sg13g2_decap_8
XFILLER_0_562 VPWR VGND sg13g2_decap_8
XFILLER_48_555 VPWR VGND sg13g2_decap_8
XFILLER_16_430 VPWR VGND sg13g2_fill_2
XFILLER_17_942 VPWR VGND sg13g2_decap_8
XFILLER_32_923 VPWR VGND sg13g2_decap_8
X_4769__64 VPWR VGND net64 sg13g2_tiehi
X_2840_ _0699_ _0762_ _0771_ VPWR VGND sg13g2_nor2_2
X_4784__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_31_466 VPWR VGND sg13g2_fill_2
X_2771_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\] _0754_ _0473_
+ VPWR VGND sg13g2_mux2_1
X_4510_ net674 net726 _0063_ VPWR VGND sg13g2_nor2_1
X_4441_ _2130_ tmds_blue.dc_balancing_reg\[4\] _2129_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_684 VPWR VGND sg13g2_decap_8
X_4372_ VPWR VGND net603 _2030_ _2064_ _2043_ _2066_ _2056_ sg13g2_a221oi_1
X_3323_ VGND VPWR _1053_ _1052_ _1046_ sg13g2_or2_1
Xfanout608 videogen.fancy_shader.video_y\[1\] net608 VPWR VGND sg13g2_buf_8
Xfanout619 net620 net619 VPWR VGND sg13g2_buf_8
X_3254_ net747 _0990_ _0991_ _0363_ VPWR VGND sg13g2_nor3_1
X_3185_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\] _0946_ _0947_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_35_750 VPWR VGND sg13g2_decap_8
XFILLER_23_934 VPWR VGND sg13g2_decap_8
XFILLER_22_477 VPWR VGND sg13g2_fill_2
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
X_2969_ videogen.fancy_shader.video_y\[5\] _0660_ _0815_ _0816_ _0817_ VPWR VGND sg13g2_nor4_1
X_4893__210 VPWR VGND net210 sg13g2_tiehi
X_4708_ net653 net704 _0259_ VPWR VGND sg13g2_nor2_1
X_4639_ net667 net718 _0192_ VPWR VGND sg13g2_nor2_1
X_4930__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_40_1026 VPWR VGND sg13g2_fill_2
XFILLER_40_252 VPWR VGND sg13g2_fill_1
XFILLER_14_978 VPWR VGND sg13g2_decap_8
XFILLER_40_263 VPWR VGND sg13g2_fill_2
XFILLER_5_665 VPWR VGND sg13g2_decap_8
XFILLER_1_860 VPWR VGND sg13g2_decap_8
XFILLER_48_330 VPWR VGND sg13g2_decap_8
XFILLER_49_897 VPWR VGND sg13g2_decap_8
X_5007__167 VPWR VGND net167 sg13g2_tiehi
X_4990_ net234 VGND VPWR _0537_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\]
+ _0185_ sg13g2_dfrbpq_1
X_3941_ _1653_ _1655_ _1667_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
X_3872_ net627 videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\]
+ net624 _1601_ VPWR VGND sg13g2_mux4_1
XFILLER_31_252 VPWR VGND sg13g2_decap_8
X_2823_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\] net778 _0767_ _0434_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_786 VPWR VGND sg13g2_decap_8
XFILLER_31_296 VPWR VGND sg13g2_fill_2
X_2754_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\] _0750_ _0486_
+ VPWR VGND sg13g2_mux2_1
X_2685_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\] net786 _0736_ _0550_
+ VPWR VGND sg13g2_mux2_1
X_4424_ _2092_ VPWR _2114_ VGND _2082_ _2090_ sg13g2_o21ai_1
X_4355_ _2018_ _2029_ _2049_ _2050_ VPWR VGND sg13g2_nor3_1
X_3306_ _1036_ _1034_ _1035_ VPWR VGND sg13g2_nand2_2
X_4286_ _0644_ _1988_ tmds_blue.n193 _1990_ VPWR VGND sg13g2_nand3_1
X_3237_ _0978_ _0979_ _0897_ _0980_ VPWR VGND sg13g2_nand3_1
X_3168_ VGND VPWR net628 _0933_ _0936_ net625 sg13g2_a21oi_1
XFILLER_27_558 VPWR VGND sg13g2_fill_2
XFILLER_14_219 VPWR VGND sg13g2_decap_8
X_3099_ VGND VPWR _0888_ _0889_ _0880_ tmds_red.dc_balancing_reg\[4\] sg13g2_a21oi_2
XFILLER_23_764 VPWR VGND sg13g2_fill_1
XFILLER_22_274 VPWR VGND sg13g2_decap_8
XFILLER_7_919 VPWR VGND sg13g2_decap_8
XFILLER_10_458 VPWR VGND sg13g2_fill_1
XFILLER_2_624 VPWR VGND sg13g2_fill_1
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_1_167 VPWR VGND sg13g2_fill_2
XFILLER_1_156 VPWR VGND sg13g2_decap_4
XFILLER_49_127 VPWR VGND sg13g2_decap_8
XFILLER_18_503 VPWR VGND sg13g2_fill_2
XFILLER_18_558 VPWR VGND sg13g2_decap_8
XFILLER_45_388 VPWR VGND sg13g2_decap_8
XFILLER_45_366 VPWR VGND sg13g2_decap_8
XFILLER_14_764 VPWR VGND sg13g2_fill_1
XFILLER_41_583 VPWR VGND sg13g2_fill_1
XFILLER_9_201 VPWR VGND sg13g2_fill_2
XFILLER_13_263 VPWR VGND sg13g2_fill_1
XFILLER_13_274 VPWR VGND sg13g2_decap_8
XFILLER_6_963 VPWR VGND sg13g2_decap_8
XFILLER_5_440 VPWR VGND sg13g2_fill_1
XFILLER_5_495 VPWR VGND sg13g2_decap_8
X_4140_ _1840_ _1854_ _1861_ _1863_ VPWR VGND sg13g2_or3_1
X_4071_ _1793_ VPWR _1794_ VGND _1778_ _1789_ sg13g2_o21ai_1
X_3022_ net439 green_tmds_par\[7\] net699 serialize.n428\[7\] VPWR VGND sg13g2_mux2_1
XFILLER_37_878 VPWR VGND sg13g2_fill_1
XFILLER_24_506 VPWR VGND sg13g2_decap_8
X_4973_ net304 VGND VPWR _0520_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\]
+ _0168_ sg13g2_dfrbpq_1
X_3924_ _1647_ _1649_ _1650_ VPWR VGND sg13g2_nor2_1
XFILLER_32_583 VPWR VGND sg13g2_decap_8
X_3855_ _1582_ _1583_ net594 _1584_ VPWR VGND sg13g2_mux2_1
X_2806_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\] _0764_ _0448_
+ VPWR VGND sg13g2_mux2_1
X_3786_ net596 VPWR _1516_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\]
+ net583 sg13g2_o21ai_1
XFILLER_30_1014 VPWR VGND sg13g2_decap_8
X_2737_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\] _0747_ _0509_
+ VPWR VGND sg13g2_mux2_1
X_2668_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\] _0733_ _0564_
+ VPWR VGND sg13g2_mux2_1
X_4407_ VPWR VGND _1989_ _2095_ _2096_ _2004_ _2098_ _2088_ sg13g2_a221oi_1
X_2599_ _0680_ _0705_ _0706_ VPWR VGND sg13g2_nor2_2
X_4338_ _2033_ _2029_ _2034_ VPWR VGND sg13g2_nor2b_1
X_4269_ _0879_ _0883_ _1974_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_823 VPWR VGND sg13g2_fill_1
XFILLER_27_344 VPWR VGND sg13g2_fill_2
XFILLER_28_845 VPWR VGND sg13g2_decap_8
XFILLER_43_826 VPWR VGND sg13g2_fill_2
XFILLER_27_377 VPWR VGND sg13g2_fill_2
X_5076__63 VPWR VGND net63 sg13g2_tiehi
XFILLER_27_399 VPWR VGND sg13g2_fill_2
XFILLER_42_347 VPWR VGND sg13g2_decap_8
XFILLER_7_716 VPWR VGND sg13g2_decap_8
XFILLER_11_778 VPWR VGND sg13g2_decap_8
XFILLER_3_911 VPWR VGND sg13g2_decap_8
XFILLER_3_988 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
Xfanout780 net781 net780 VPWR VGND sg13g2_buf_8
XFILLER_18_344 VPWR VGND sg13g2_decap_8
XFILLER_45_163 VPWR VGND sg13g2_fill_2
XFILLER_18_388 VPWR VGND sg13g2_fill_2
X_5043__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_33_347 VPWR VGND sg13g2_fill_2
XFILLER_14_583 VPWR VGND sg13g2_decap_4
X_3640_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\] net584 _1370_ VPWR
+ VGND sg13g2_nor2_1
X_3571_ _1300_ VPWR _1301_ VGND _1264_ _1276_ sg13g2_o21ai_1
X_2522_ VPWR _0640_ videogen.fancy_shader.video_x\[5\] VGND sg13g2_inv_1
X_4123_ _1826_ VPWR _1846_ VGND _1806_ _1829_ sg13g2_o21ai_1
X_4054_ _1777_ _1773_ _1776_ VPWR VGND sg13g2_nand2_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_2
X_3005_ net426 blue_tmds_par\[1\] net699 serialize.n429\[1\] VPWR VGND sg13g2_mux2_1
XFILLER_37_653 VPWR VGND sg13g2_decap_8
X_4956_ net389 VGND VPWR _0503_ tmds_red.dc_balancing_reg\[2\] net647 sg13g2_dfrbpq_2
X_4887_ net222 VGND VPWR _0438_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\]
+ _0095_ sg13g2_dfrbpq_1
X_3907_ _1633_ _1063_ _1631_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_380 VPWR VGND sg13g2_decap_8
X_3838_ _1567_ _0674_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
X_3769_ _1498_ VPWR _1499_ VGND _1462_ _1474_ sg13g2_o21ai_1
XFILLER_10_23 VPWR VGND sg13g2_decap_8
XFILLER_0_947 VPWR VGND sg13g2_decap_8
X_4712__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_19_10 VPWR VGND sg13g2_decap_8
XFILLER_19_108 VPWR VGND sg13g2_fill_2
XFILLER_27_185 VPWR VGND sg13g2_decap_8
XFILLER_28_686 VPWR VGND sg13g2_fill_2
XFILLER_15_347 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_fill_2
XFILLER_31_818 VPWR VGND sg13g2_decap_8
XFILLER_11_531 VPWR VGND sg13g2_fill_1
XFILLER_7_535 VPWR VGND sg13g2_fill_1
XFILLER_3_730 VPWR VGND sg13g2_fill_2
XFILLER_19_631 VPWR VGND sg13g2_fill_1
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_19_675 VPWR VGND sg13g2_decap_8
XFILLER_34_623 VPWR VGND sg13g2_fill_1
X_4810_ net354 VGND VPWR _0361_ videogen.fancy_shader.video_y\[5\] net636 sg13g2_dfrbpq_2
X_4948__37 VPWR VGND net37 sg13g2_tiehi
XFILLER_21_306 VPWR VGND sg13g2_decap_8
XFILLER_34_689 VPWR VGND sg13g2_decap_8
X_4741_ net109 VGND VPWR _0292_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\]
+ _0023_ sg13g2_dfrbpq_1
X_4672_ net671 net722 _0225_ VPWR VGND sg13g2_nor2_1
X_3623_ net618 VPWR _1353_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\]
+ net575 sg13g2_o21ai_1
XFILLER_30_895 VPWR VGND sg13g2_decap_8
X_3554_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\] net563 _1284_ VPWR
+ VGND sg13g2_nor2_1
X_3485_ _1215_ _1212_ _1214_ VPWR VGND sg13g2_nand2_1
X_5086_ net799 VGND VPWR serialize.n428\[1\] serialize.n455 clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4106_ VGND VPWR _1827_ _1828_ _1829_ _1823_ sg13g2_a21oi_1
X_4926__120 VPWR VGND net120 sg13g2_tiehi
X_4037_ _1760_ _1755_ _1759_ VPWR VGND sg13g2_nand2_1
XFILLER_12_306 VPWR VGND sg13g2_fill_2
XFILLER_24_188 VPWR VGND sg13g2_decap_8
X_4939_ net74 VGND VPWR _0486_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\]
+ _0143_ sg13g2_dfrbpq_1
XFILLER_21_884 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_0_744 VPWR VGND sg13g2_decap_8
XFILLER_46_74 VPWR VGND sg13g2_fill_2
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_29_995 VPWR VGND sg13g2_decap_8
XFILLER_15_177 VPWR VGND sg13g2_decap_8
XFILLER_30_136 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_12_873 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_8_877 VPWR VGND sg13g2_decap_8
X_3270_ _1001_ _0667_ _1000_ VPWR VGND sg13g2_nand2_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_35_921 VPWR VGND sg13g2_fill_2
XFILLER_22_626 VPWR VGND sg13g2_decap_8
XFILLER_35_998 VPWR VGND sg13g2_decap_8
X_2985_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0825_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\]
+ _0829_ VPWR VGND sg13g2_nand3_1
X_4724_ net139 VGND VPWR _0275_ red_tmds_par\[1\] net647 sg13g2_dfrbpq_1
X_4655_ net669 net719 _0208_ VPWR VGND sg13g2_nor2_1
X_4586_ net677 net729 _0139_ VPWR VGND sg13g2_nor2_1
X_3606_ net623 VPWR _1336_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\]
+ net562 sg13g2_o21ai_1
X_3537_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\] net564 _1267_ VPWR
+ VGND sg13g2_nor2_1
X_3468_ VGND VPWR _1112_ _1121_ _1198_ _1124_ sg13g2_a21oi_1
X_3399_ _1120_ _1124_ _1129_ VPWR VGND sg13g2_nor2_1
XFILLER_29_236 VPWR VGND sg13g2_decap_8
XFILLER_45_718 VPWR VGND sg13g2_decap_8
XFILLER_44_206 VPWR VGND sg13g2_fill_2
XFILLER_38_792 VPWR VGND sg13g2_fill_1
X_5069_ net177 VGND VPWR _0616_ blue_tmds_par\[7\] net642 sg13g2_dfrbpq_1
XFILLER_37_280 VPWR VGND sg13g2_fill_1
XFILLER_25_420 VPWR VGND sg13g2_fill_1
XFILLER_26_954 VPWR VGND sg13g2_decap_8
XFILLER_13_626 VPWR VGND sg13g2_fill_2
XFILLER_16_55 VPWR VGND sg13g2_fill_1
XFILLER_12_103 VPWR VGND sg13g2_fill_1
XFILLER_12_114 VPWR VGND sg13g2_decap_8
XFILLER_41_979 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_40_489 VPWR VGND sg13g2_fill_1
X_5000__195 VPWR VGND net195 sg13g2_tiehi
XFILLER_5_825 VPWR VGND sg13g2_decap_4
XFILLER_0_541 VPWR VGND sg13g2_decap_8
XFILLER_48_534 VPWR VGND sg13g2_decap_8
XFILLER_36_707 VPWR VGND sg13g2_fill_1
XFILLER_17_921 VPWR VGND sg13g2_decap_8
X_4842__313 VPWR VGND net313 sg13g2_tiehi
XFILLER_17_998 VPWR VGND sg13g2_decap_8
XFILLER_32_902 VPWR VGND sg13g2_decap_8
X_2770_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\] _0754_ _0474_
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_681 VPWR VGND sg13g2_decap_8
XFILLER_11_191 VPWR VGND sg13g2_fill_2
X_4440_ _2128_ VPWR _2129_ VGND tmds_blue.dc_balancing_reg\[3\] _2080_ sg13g2_o21ai_1
X_4941__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_4_880 VPWR VGND sg13g2_decap_8
X_4371_ _2031_ _2058_ net602 _2065_ VPWR VGND _2064_ sg13g2_nand4_1
X_3322_ _1051_ _1049_ _1052_ VPWR VGND sg13g2_xor2_1
Xfanout609 videogen.fancy_shader.video_y\[0\] net609 VPWR VGND sg13g2_buf_8
X_3253_ _0991_ videogen.fancy_shader.video_y\[7\] videogen.fancy_shader.video_y\[6\]
+ _0988_ VPWR VGND sg13g2_and3_1
XFILLER_39_534 VPWR VGND sg13g2_decap_8
X_3184_ _0944_ _0945_ _0946_ _0330_ VPWR VGND sg13g2_nor3_1
XFILLER_23_913 VPWR VGND sg13g2_decap_8
X_2968_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\] videogen.fancy_shader.video_y\[4\]
+ _0816_ VPWR VGND sg13g2_nand3_1
XFILLER_31_990 VPWR VGND sg13g2_decap_8
X_4707_ net654 net705 _0258_ VPWR VGND sg13g2_nor2_1
X_4638_ net666 net717 _0191_ VPWR VGND sg13g2_nor2_1
X_2899_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\] _0784_ _0301_
+ VPWR VGND sg13g2_mux2_1
XFILLER_2_839 VPWR VGND sg13g2_decap_8
X_4569_ net676 net728 _0122_ VPWR VGND sg13g2_nor2_1
XFILLER_1_349 VPWR VGND sg13g2_fill_1
XFILLER_40_1005 VPWR VGND sg13g2_decap_8
XFILLER_17_206 VPWR VGND sg13g2_decap_8
XFILLER_26_773 VPWR VGND sg13g2_decap_4
XFILLER_41_732 VPWR VGND sg13g2_fill_1
XFILLER_40_220 VPWR VGND sg13g2_decap_8
XFILLER_14_957 VPWR VGND sg13g2_decap_8
XFILLER_25_261 VPWR VGND sg13g2_fill_1
XFILLER_25_294 VPWR VGND sg13g2_fill_1
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_9_405 VPWR VGND sg13g2_decap_8
XFILLER_40_275 VPWR VGND sg13g2_fill_1
XFILLER_13_489 VPWR VGND sg13g2_fill_2
XFILLER_5_699 VPWR VGND sg13g2_fill_2
XFILLER_4_176 VPWR VGND sg13g2_fill_1
XFILLER_49_876 VPWR VGND sg13g2_decap_8
XFILLER_48_386 VPWR VGND sg13g2_decap_8
X_5046__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_1_1021 VPWR VGND sg13g2_decap_8
XFILLER_36_537 VPWR VGND sg13g2_decap_8
X_3940_ _1666_ _1663_ _1664_ _1661_ _1657_ VPWR VGND sg13g2_a22oi_1
XFILLER_17_751 VPWR VGND sg13g2_fill_2
XFILLER_44_592 VPWR VGND sg13g2_decap_8
XFILLER_16_272 VPWR VGND sg13g2_decap_8
X_3871_ net624 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\]
+ net627 _1600_ VPWR VGND sg13g2_mux4_1
XFILLER_32_765 VPWR VGND sg13g2_decap_8
X_2822_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\] net767 _0767_ _0435_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_949 VPWR VGND sg13g2_decap_8
XFILLER_31_275 VPWR VGND sg13g2_decap_4
X_2753_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\] _0750_ _0487_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
X_2684_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\] net775 _0736_ _0551_
+ VPWR VGND sg13g2_mux2_1
X_4423_ _2113_ _2104_ _2111_ VPWR VGND sg13g2_xnor2_1
X_4354_ _2047_ _2046_ _2049_ VPWR VGND sg13g2_xor2_1
X_3305_ _1035_ net546 _1027_ VPWR VGND sg13g2_nand2b_1
X_4285_ _1989_ _0644_ VPWR VGND _1988_ sg13g2_nand2b_2
XFILLER_39_342 VPWR VGND sg13g2_fill_1
X_3236_ _0632_ videogen.fancy_shader.video_y\[8\] _0815_ _0911_ _0979_ VPWR VGND sg13g2_nor4_1
X_3167_ net578 _0931_ _0932_ _0935_ VPWR VGND sg13g2_nor3_1
XFILLER_27_537 VPWR VGND sg13g2_fill_2
X_3098_ tmds_red.dc_balancing_reg\[4\] _0856_ _0887_ _0888_ VPWR VGND sg13g2_nor3_1
XFILLER_35_570 VPWR VGND sg13g2_decap_8
XFILLER_10_426 VPWR VGND sg13g2_fill_1
XFILLER_11_949 VPWR VGND sg13g2_decap_8
XFILLER_22_264 VPWR VGND sg13g2_decap_4
XFILLER_23_798 VPWR VGND sg13g2_decap_8
X_4771__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_38_53 VPWR VGND sg13g2_decap_4
XFILLER_38_42 VPWR VGND sg13g2_fill_1
XFILLER_46_846 VPWR VGND sg13g2_fill_2
XFILLER_46_879 VPWR VGND sg13g2_decap_8
XFILLER_14_721 VPWR VGND sg13g2_decap_4
X_4906__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_9_235 VPWR VGND sg13g2_fill_2
XFILLER_10_982 VPWR VGND sg13g2_decap_8
XFILLER_6_942 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
XFILLER_49_651 VPWR VGND sg13g2_fill_1
X_4070_ net547 _1234_ _1793_ VPWR VGND sg13g2_nor2_1
XFILLER_23_1011 VPWR VGND sg13g2_decap_8
X_3021_ net427 green_tmds_par\[6\] net696 serialize.n428\[6\] VPWR VGND sg13g2_mux2_1
XFILLER_37_857 VPWR VGND sg13g2_decap_4
XFILLER_36_323 VPWR VGND sg13g2_decap_4
X_4972_ net308 VGND VPWR _0519_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\]
+ _0167_ sg13g2_dfrbpq_1
X_3923_ _1640_ _1641_ _1649_ VPWR VGND sg13g2_and2_1
X_3854_ net626 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\]
+ net625 _1583_ VPWR VGND sg13g2_mux4_1
X_2805_ _0764_ _0710_ _0763_ VPWR VGND sg13g2_nand2_2
X_3785_ _1511_ _1512_ _1513_ _1514_ _1515_ VPWR VGND sg13g2_nor4_1
X_2736_ _0747_ _0702_ _0720_ VPWR VGND sg13g2_nand2_2
X_2667_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\] _0733_ _0565_
+ VPWR VGND sg13g2_mux2_1
X_4406_ VPWR _2097_ _2096_ VGND sg13g2_inv_1
X_2598_ _0682_ _0685_ net543 _0705_ VPWR VGND sg13g2_nand3_1
X_4337_ _0841_ VPWR _2033_ VGND tmds_green.dc_balancing_reg\[1\] _0842_ sg13g2_o21ai_1
X_4268_ VGND VPWR _1955_ _1956_ _1973_ _1958_ sg13g2_a21oi_1
X_3219_ _0968_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.n646\[5\] _0965_
+ VPWR VGND sg13g2_and3_1
X_4199_ net803 _1915_ _0385_ VPWR VGND sg13g2_and2_1
XFILLER_15_518 VPWR VGND sg13g2_fill_1
XFILLER_28_879 VPWR VGND sg13g2_decap_8
XFILLER_42_359 VPWR VGND sg13g2_fill_1
XFILLER_11_702 VPWR VGND sg13g2_decap_8
XFILLER_23_562 VPWR VGND sg13g2_decap_8
XFILLER_10_234 VPWR VGND sg13g2_fill_1
XFILLER_6_227 VPWR VGND sg13g2_decap_4
XFILLER_40_87 VPWR VGND sg13g2_fill_2
XFILLER_40_76 VPWR VGND sg13g2_decap_8
XFILLER_3_967 VPWR VGND sg13g2_decap_8
XFILLER_2_433 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_2_488 VPWR VGND sg13g2_decap_8
Xfanout770 net771 net770 VPWR VGND sg13g2_buf_8
Xfanout792 ui_in[4] net792 VPWR VGND sg13g2_buf_8
XFILLER_18_301 VPWR VGND sg13g2_decap_4
XFILLER_19_824 VPWR VGND sg13g2_fill_1
Xfanout781 ui_in[5] net781 VPWR VGND sg13g2_buf_8
XFILLER_19_879 VPWR VGND sg13g2_decap_8
XFILLER_46_698 VPWR VGND sg13g2_fill_2
X_3570_ _0636_ _1299_ _1300_ VPWR VGND sg13g2_nor2_1
X_5050__114 VPWR VGND net114 sg13g2_tiehi
X_2521_ VPWR _0639_ net619 VGND sg13g2_inv_1
X_4122_ _1845_ _1839_ _1844_ VPWR VGND sg13g2_nand2_1
X_4053_ _1774_ VPWR _1776_ VGND _1765_ _1775_ sg13g2_o21ai_1
X_3004_ net433 blue_tmds_par\[0\] net699 serialize.n429\[0\] VPWR VGND sg13g2_mux2_1
XFILLER_25_816 VPWR VGND sg13g2_decap_8
XFILLER_36_142 VPWR VGND sg13g2_fill_2
XFILLER_18_890 VPWR VGND sg13g2_decap_4
XFILLER_25_849 VPWR VGND sg13g2_fill_1
XFILLER_36_164 VPWR VGND sg13g2_decap_4
X_4955_ net391 VGND VPWR _0502_ tmds_red.dc_balancing_reg\[1\] net647 sg13g2_dfrbpq_2
X_3906_ net546 _1052_ _1063_ _1626_ _1632_ VPWR VGND sg13g2_and4_1
X_4886_ net224 VGND VPWR _0437_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\]
+ _0094_ sg13g2_dfrbpq_1
XFILLER_20_521 VPWR VGND sg13g2_decap_8
X_3837_ VGND VPWR _1566_ net573 videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\]
+ sg13g2_or2_1
XFILLER_20_587 VPWR VGND sg13g2_decap_4
X_3768_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1497_ _1498_ VPWR VGND
+ sg13g2_nor2_1
X_2719_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\] _0743_ _0523_
+ VPWR VGND sg13g2_mux2_1
X_3699_ net616 VPWR _1429_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\]
+ net578 sg13g2_o21ai_1
XFILLER_0_926 VPWR VGND sg13g2_decap_8
XFILLER_47_407 VPWR VGND sg13g2_fill_2
XFILLER_16_816 VPWR VGND sg13g2_decap_8
XFILLER_27_153 VPWR VGND sg13g2_decap_8
XFILLER_43_613 VPWR VGND sg13g2_fill_1
XFILLER_42_156 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_4
XFILLER_11_510 VPWR VGND sg13g2_decap_8
XFILLER_7_503 VPWR VGND sg13g2_fill_2
XFILLER_13_1021 VPWR VGND sg13g2_decap_8
XFILLER_39_919 VPWR VGND sg13g2_decap_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_19_654 VPWR VGND sg13g2_fill_1
XFILLER_46_495 VPWR VGND sg13g2_fill_1
X_4880__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_33_178 VPWR VGND sg13g2_fill_1
X_4740_ net111 VGND VPWR _0291_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\]
+ _0022_ sg13g2_dfrbpq_1
XFILLER_33_189 VPWR VGND sg13g2_fill_2
X_4671_ net686 net737 _0224_ VPWR VGND sg13g2_nor2_1
XFILLER_30_852 VPWR VGND sg13g2_decap_8
XFILLER_30_863 VPWR VGND sg13g2_fill_2
XFILLER_30_874 VPWR VGND sg13g2_decap_8
X_3622_ _1351_ _1352_ VPWR VGND sg13g2_inv_4
X_3553_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\] net553 _1283_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_44_0 VPWR VGND sg13g2_decap_4
X_3484_ _1214_ net544 _1209_ VPWR VGND sg13g2_nand2_1
X_4105_ _1811_ _1822_ _1828_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_418 VPWR VGND sg13g2_fill_1
X_5085_ net799 VGND VPWR serialize.n428\[0\] serialize.n453 clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4036_ _1744_ VPWR _1759_ VGND _1735_ _1748_ sg13g2_o21ai_1
XFILLER_25_635 VPWR VGND sg13g2_decap_8
XFILLER_13_819 VPWR VGND sg13g2_decap_4
XFILLER_25_679 VPWR VGND sg13g2_decap_8
X_4938_ net88 VGND VPWR _0485_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\]
+ _0142_ sg13g2_dfrbpq_1
X_4869_ net261 VGND VPWR _0420_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\]
+ _0077_ sg13g2_dfrbpq_1
XFILLER_4_506 VPWR VGND sg13g2_decap_8
XFILLER_21_89 VPWR VGND sg13g2_decap_4
XFILLER_0_723 VPWR VGND sg13g2_decap_8
XFILLER_48_705 VPWR VGND sg13g2_fill_2
XFILLER_29_974 VPWR VGND sg13g2_decap_8
XFILLER_46_64 VPWR VGND sg13g2_fill_2
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_4
XFILLER_28_495 VPWR VGND sg13g2_fill_2
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_43_498 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_fill_1
XFILLER_38_204 VPWR VGND sg13g2_fill_2
X_2984_ VGND VPWR _0818_ _0828_ net19 _0820_ sg13g2_a21oi_1
XFILLER_21_126 VPWR VGND sg13g2_decap_4
XFILLER_34_487 VPWR VGND sg13g2_decap_4
X_4723_ net140 VGND VPWR _0274_ red_tmds_par\[0\] net647 sg13g2_dfrbpq_1
X_4654_ net684 net719 _0207_ VPWR VGND sg13g2_nor2_1
X_4585_ net676 net728 _0138_ VPWR VGND sg13g2_nor2_1
X_3605_ net599 _1329_ _1334_ _1335_ VPWR VGND sg13g2_nor3_1
X_3536_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\] net577 _1266_ VPWR
+ VGND sg13g2_nor2_1
X_3467_ _1066_ _1192_ _1193_ _1196_ _1197_ VPWR VGND sg13g2_or4_1
X_3398_ _1113_ _1120_ _1066_ _1128_ VPWR VGND _1126_ sg13g2_nand4_1
X_5068_ net185 VGND VPWR _0615_ blue_tmds_par\[6\] net642 sg13g2_dfrbpq_1
X_4019_ VPWR _1742_ _1741_ VGND sg13g2_inv_1
XFILLER_26_933 VPWR VGND sg13g2_decap_8
XFILLER_41_958 VPWR VGND sg13g2_decap_8
XFILLER_13_649 VPWR VGND sg13g2_decap_8
XFILLER_32_66 VPWR VGND sg13g2_decap_4
XFILLER_4_303 VPWR VGND sg13g2_fill_2
XFILLER_10_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_597 VPWR VGND sg13g2_decap_8
XFILLER_16_421 VPWR VGND sg13g2_fill_1
XFILLER_16_432 VPWR VGND sg13g2_fill_1
XFILLER_44_763 VPWR VGND sg13g2_fill_2
XFILLER_43_240 VPWR VGND sg13g2_fill_1
XFILLER_16_443 VPWR VGND sg13g2_fill_1
XFILLER_16_454 VPWR VGND sg13g2_fill_2
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_43_284 VPWR VGND sg13g2_fill_2
XFILLER_31_435 VPWR VGND sg13g2_fill_2
XFILLER_32_969 VPWR VGND sg13g2_decap_8
XFILLER_40_991 VPWR VGND sg13g2_decap_8
XFILLER_8_664 VPWR VGND sg13g2_decap_8
XFILLER_7_163 VPWR VGND sg13g2_decap_8
X_4916__164 VPWR VGND net164 sg13g2_tiehi
X_4370_ _2064_ _2015_ _2029_ VPWR VGND sg13g2_nand2b_1
X_3321_ _1051_ videogen.fancy_shader.video_y\[4\] videogen.fancy_shader.n646\[4\]
+ VPWR VGND sg13g2_xnor2_1
X_4732__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_3_391 VPWR VGND sg13g2_decap_8
X_3252_ VGND VPWR videogen.fancy_shader.video_y\[6\] _0988_ _0990_ videogen.fancy_shader.video_y\[7\]
+ sg13g2_a21oi_1
X_3183_ _0914_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0946_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_27_708 VPWR VGND sg13g2_decap_8
XFILLER_34_240 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_fill_1
XFILLER_23_969 VPWR VGND sg13g2_decap_8
X_2967_ _0815_ net608 net609 VPWR VGND sg13g2_nand2_1
X_2898_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\] _0784_ _0302_
+ VPWR VGND sg13g2_mux2_1
X_4706_ _1994_ _1998_ _0614_ VPWR VGND sg13g2_nor2_1
X_4637_ net667 net717 _0190_ VPWR VGND sg13g2_nor2_1
XFILLER_2_818 VPWR VGND sg13g2_decap_8
X_4568_ net681 net734 _0121_ VPWR VGND sg13g2_nor2_1
X_4499_ net652 net703 _0052_ VPWR VGND sg13g2_nor2_1
X_3519_ _1246_ _1234_ _1247_ _1249_ VPWR VGND sg13g2_a21o_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_11 VPWR VGND sg13g2_decap_4
XFILLER_14_936 VPWR VGND sg13g2_decap_8
XFILLER_25_273 VPWR VGND sg13g2_decap_8
XFILLER_43_54 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_22_991 VPWR VGND sg13g2_decap_8
X_4766__69 VPWR VGND net69 sg13g2_tiehi
X_4952__397 VPWR VGND net397 sg13g2_tiehi
XFILLER_4_188 VPWR VGND sg13g2_decap_8
XFILLER_0_372 VPWR VGND sg13g2_fill_2
XFILLER_1_895 VPWR VGND sg13g2_decap_8
XFILLER_49_855 VPWR VGND sg13g2_decap_8
XFILLER_48_365 VPWR VGND sg13g2_decap_8
XFILLER_1_1000 VPWR VGND sg13g2_decap_8
XFILLER_17_796 VPWR VGND sg13g2_fill_2
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
X_3870_ _0636_ _1590_ _1598_ _1599_ VPWR VGND sg13g2_nor3_1
X_2821_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\] net757 _0767_ _0436_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_928 VPWR VGND sg13g2_decap_8
XFILLER_31_298 VPWR VGND sg13g2_fill_1
X_2752_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\] _0750_ _0488_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_4422_ _2111_ VPWR _2112_ VGND _2085_ _2087_ sg13g2_o21ai_1
X_2683_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\] net766 _0736_ _0552_
+ VPWR VGND sg13g2_mux2_1
X_4353_ VPWR _2048_ _2047_ VGND sg13g2_inv_1
X_4284_ tmds_blue.dc_balancing_reg\[0\] tmds_blue.dc_balancing_reg\[1\] tmds_blue.dc_balancing_reg\[3\]
+ tmds_blue.dc_balancing_reg\[2\] _1988_ VPWR VGND sg13g2_or4_1
X_3304_ _1034_ _1027_ net546 VPWR VGND sg13g2_nand2b_1
X_3235_ videogen.fancy_shader.video_y\[7\] videogen.fancy_shader.video_y\[6\] videogen.fancy_shader.video_y\[5\]
+ videogen.fancy_shader.video_y\[4\] _0978_ VPWR VGND sg13g2_nor4_1
X_3166_ _0793_ _0934_ _0324_ VPWR VGND sg13g2_nor2_1
X_3097_ _0878_ _0886_ _0887_ VPWR VGND sg13g2_nor2_1
XFILLER_42_519 VPWR VGND sg13g2_decap_8
XFILLER_11_928 VPWR VGND sg13g2_decap_8
XFILLER_23_777 VPWR VGND sg13g2_decap_8
X_3999_ VGND VPWR _1450_ _1451_ _1723_ _1549_ sg13g2_a21oi_1
XFILLER_6_409 VPWR VGND sg13g2_decap_8
XFILLER_1_169 VPWR VGND sg13g2_fill_1
XFILLER_46_803 VPWR VGND sg13g2_decap_8
XFILLER_18_505 VPWR VGND sg13g2_fill_1
XFILLER_33_519 VPWR VGND sg13g2_decap_8
XFILLER_26_582 VPWR VGND sg13g2_decap_8
XFILLER_41_530 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_fill_1
XFILLER_9_214 VPWR VGND sg13g2_fill_1
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_10_961 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_4987__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_49_630 VPWR VGND sg13g2_decap_8
X_3020_ _0834_ VPWR serialize.n428\[5\] VGND _0657_ net700 sg13g2_o21ai_1
XFILLER_0_191 VPWR VGND sg13g2_decap_8
X_4971_ net312 VGND VPWR _0518_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\]
+ _0166_ sg13g2_dfrbpq_1
X_3922_ _1647_ _1643_ _1648_ VPWR VGND sg13g2_xor2_1
X_3853_ net627 videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\]
+ net624 _1582_ VPWR VGND sg13g2_mux4_1
X_2804_ VPWR _0763_ _0762_ VGND sg13g2_inv_1
XFILLER_32_596 VPWR VGND sg13g2_fill_2
X_3784_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\] net549 _1514_ VPWR
+ VGND sg13g2_nor2_1
X_2735_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\] _0746_ _0510_
+ VPWR VGND sg13g2_mux2_1
X_2666_ _0733_ _0715_ _0731_ VPWR VGND sg13g2_nand2_2
X_4405_ _2091_ _2093_ _2096_ VPWR VGND sg13g2_nor2b_1
X_5031__295 VPWR VGND net295 sg13g2_tiehi
X_2597_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\] _0704_ _0606_
+ VPWR VGND sg13g2_mux2_1
X_4336_ _2029_ _2016_ _2032_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
X_4267_ net570 _1972_ _0504_ VPWR VGND sg13g2_nor2_1
X_3218_ VGND VPWR videogen.fancy_shader.n646\[5\] _0965_ _0967_ videogen.fancy_shader.n646\[6\]
+ sg13g2_a21oi_1
X_4198_ _1914_ VPWR _1915_ VGND _0891_ _1913_ sg13g2_o21ai_1
X_3149_ _0919_ _0921_ _0922_ _0319_ VPWR VGND sg13g2_nor3_1
XFILLER_27_313 VPWR VGND sg13g2_decap_4
XFILLER_27_346 VPWR VGND sg13g2_fill_1
XFILLER_27_357 VPWR VGND sg13g2_fill_2
XFILLER_43_839 VPWR VGND sg13g2_decap_4
XFILLER_27_379 VPWR VGND sg13g2_fill_1
XFILLER_23_541 VPWR VGND sg13g2_decap_8
XFILLER_35_390 VPWR VGND sg13g2_decap_4
XFILLER_24_45 VPWR VGND sg13g2_decap_4
XFILLER_11_758 VPWR VGND sg13g2_decap_4
XFILLER_3_946 VPWR VGND sg13g2_decap_8
XFILLER_46_1012 VPWR VGND sg13g2_decap_8
X_5084__403 VPWR VGND net403 sg13g2_tiehi
XFILLER_49_42 VPWR VGND sg13g2_decap_8
Xfanout760 net761 net760 VPWR VGND sg13g2_buf_8
Xfanout771 ui_in[6] net771 VPWR VGND sg13g2_buf_8
Xfanout793 net794 net793 VPWR VGND sg13g2_buf_8
Xfanout782 net792 net782 VPWR VGND sg13g2_buf_8
XFILLER_46_622 VPWR VGND sg13g2_fill_1
XFILLER_19_847 VPWR VGND sg13g2_decap_8
XFILLER_46_655 VPWR VGND sg13g2_decap_4
XFILLER_45_165 VPWR VGND sg13g2_fill_1
XFILLER_27_891 VPWR VGND sg13g2_decap_8
XFILLER_33_327 VPWR VGND sg13g2_decap_8
XFILLER_33_349 VPWR VGND sg13g2_fill_1
XFILLER_41_393 VPWR VGND sg13g2_fill_2
XFILLER_41_371 VPWR VGND sg13g2_decap_8
X_4839__319 VPWR VGND net319 sg13g2_tiehi
XFILLER_10_791 VPWR VGND sg13g2_fill_2
X_2520_ VPWR _0638_ net614 VGND sg13g2_inv_1
XFILLER_6_795 VPWR VGND sg13g2_decap_4
X_4121_ _1830_ _1842_ _1844_ VPWR VGND sg13g2_nor2_1
X_4850__298 VPWR VGND net298 sg13g2_tiehi
X_4052_ _1775_ _1767_ _1762_ _1764_ _1758_ VPWR VGND sg13g2_a22oi_1
X_3003_ VGND VPWR serialize.n431\[6\] serialize.n410 net415 sg13g2_or2_1
XFILLER_37_611 VPWR VGND sg13g2_decap_8
XFILLER_37_699 VPWR VGND sg13g2_decap_8
X_4954_ net393 VGND VPWR _0501_ tmds_red.dc_balancing_reg\[0\] net647 sg13g2_dfrbpq_1
X_3905_ _1052_ _1626_ net546 _1631_ VPWR VGND sg13g2_nand3_1
X_4885_ net226 VGND VPWR _0436_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\]
+ _0093_ sg13g2_dfrbpq_1
X_3836_ VGND VPWR _1565_ net561 videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\]
+ sg13g2_or2_1
XFILLER_20_566 VPWR VGND sg13g2_decap_8
X_3767_ net612 _1485_ _1496_ _1497_ VPWR VGND sg13g2_nor3_1
X_2718_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\] _0743_ _0524_
+ VPWR VGND sg13g2_mux2_1
X_3698_ _1424_ _1425_ _1426_ _1427_ _1428_ VPWR VGND sg13g2_nor4_1
XFILLER_10_58 VPWR VGND sg13g2_decap_4
XFILLER_0_905 VPWR VGND sg13g2_decap_8
X_2649_ net600 _0673_ net626 _0728_ VPWR VGND _0696_ sg13g2_nand4_1
XFILLER_48_909 VPWR VGND sg13g2_decap_8
X_4319_ _2016_ net601 VPWR VGND tmds_green.dc_balancing_reg\[1\] sg13g2_nand2b_2
XFILLER_47_419 VPWR VGND sg13g2_fill_2
XFILLER_28_633 VPWR VGND sg13g2_decap_4
XFILLER_27_143 VPWR VGND sg13g2_decap_4
XFILLER_28_699 VPWR VGND sg13g2_decap_4
X_5003__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_42_168 VPWR VGND sg13g2_fill_2
XFILLER_24_883 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_fill_2
X_4977__289 VPWR VGND net289 sg13g2_tiehi
XFILLER_13_1000 VPWR VGND sg13g2_decap_8
XFILLER_3_798 VPWR VGND sg13g2_decap_8
XFILLER_2_253 VPWR VGND sg13g2_fill_1
XFILLER_38_408 VPWR VGND sg13g2_decap_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_18_8 VPWR VGND sg13g2_decap_8
Xfanout590 net591 net590 VPWR VGND sg13g2_buf_8
XFILLER_18_110 VPWR VGND sg13g2_decap_8
XFILLER_18_132 VPWR VGND sg13g2_fill_2
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_33_135 VPWR VGND sg13g2_fill_1
X_4670_ net671 net722 _0223_ VPWR VGND sg13g2_nor2_1
X_3621_ _1350_ VPWR _1351_ VGND net2 _0651_ sg13g2_o21ai_1
X_3552_ net621 VPWR _1282_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\]
+ net578 sg13g2_o21ai_1
X_3483_ VGND VPWR _1207_ _1209_ _1213_ net544 sg13g2_a21oi_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_5_1009 VPWR VGND sg13g2_decap_8
X_4104_ _1806_ _1821_ _1824_ _1825_ _1827_ VPWR VGND sg13g2_or4_1
X_5084_ net403 VGND VPWR _0631_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\]
+ _0261_ sg13g2_dfrbpq_1
X_4035_ _1749_ VPWR _1758_ VGND _1753_ _1757_ sg13g2_o21ai_1
XFILLER_38_986 VPWR VGND sg13g2_decap_8
X_4742__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
X_4937_ net92 VGND VPWR _0001_ videogen.test_lut_thingy.pixel_feeder_inst.state\[3\]
+ net634 sg13g2_dfrbpq_1
XFILLER_21_820 VPWR VGND sg13g2_decap_8
X_4868_ net263 VGND VPWR _0419_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\]
+ _0076_ sg13g2_dfrbpq_1
XFILLER_21_842 VPWR VGND sg13g2_decap_8
X_3819_ _1548_ _1451_ _1549_ VPWR VGND sg13g2_nor2b_2
X_4799_ net376 VGND VPWR _0350_ videogen.fancy_shader.n646\[4\] net637 sg13g2_dfrbpq_2
XFILLER_0_702 VPWR VGND sg13g2_decap_8
XFILLER_43_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_779 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_fill_2
XFILLER_29_953 VPWR VGND sg13g2_decap_8
XFILLER_46_76 VPWR VGND sg13g2_fill_1
XFILLER_28_474 VPWR VGND sg13g2_decap_8
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_fill_1
XFILLER_15_146 VPWR VGND sg13g2_fill_2
XFILLER_15_168 VPWR VGND sg13g2_decap_4
XFILLER_30_127 VPWR VGND sg13g2_fill_2
XFILLER_7_312 VPWR VGND sg13g2_fill_2
XFILLER_4_1020 VPWR VGND sg13g2_decap_8
XFILLER_35_956 VPWR VGND sg13g2_fill_1
X_2983_ _0828_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0825_ VPWR VGND
+ sg13g2_xnor2_1
X_4722_ net141 VGND VPWR _0273_ green_tmds_par\[7\] net646 sg13g2_dfrbpq_1
XFILLER_21_149 VPWR VGND sg13g2_fill_2
X_4944__53 VPWR VGND net53 sg13g2_tiehi
X_4653_ net669 net720 _0206_ VPWR VGND sg13g2_nor2_1
X_3604_ _1330_ _1331_ _1332_ _1333_ _1334_ VPWR VGND sg13g2_nor4_1
X_4584_ net677 net729 _0137_ VPWR VGND sg13g2_nor2_1
X_3535_ net594 VPWR _1265_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\]
+ net586 sg13g2_o21ai_1
X_3466_ _1121_ VPWR _1196_ VGND net542 _1124_ sg13g2_o21ai_1
X_3397_ _1113_ _1126_ _1127_ VPWR VGND sg13g2_and2_1
X_5067_ net193 VGND VPWR _0614_ blue_tmds_par\[5\] net641 sg13g2_dfrbpq_1
XFILLER_44_219 VPWR VGND sg13g2_fill_1
X_4018_ _1737_ _1637_ _1741_ VPWR VGND sg13g2_xor2_1
XFILLER_26_912 VPWR VGND sg13g2_decap_8
XFILLER_16_35 VPWR VGND sg13g2_decap_4
XFILLER_41_926 VPWR VGND sg13g2_decap_8
XFILLER_26_989 VPWR VGND sg13g2_decap_8
XFILLER_13_628 VPWR VGND sg13g2_fill_1
XFILLER_20_160 VPWR VGND sg13g2_fill_1
XFILLER_10_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_337 VPWR VGND sg13g2_fill_2
XFILLER_48_514 VPWR VGND sg13g2_fill_2
XFILLER_0_576 VPWR VGND sg13g2_decap_8
XFILLER_48_569 VPWR VGND sg13g2_decap_8
XFILLER_29_750 VPWR VGND sg13g2_fill_2
XFILLER_29_772 VPWR VGND sg13g2_decap_4
XFILLER_17_956 VPWR VGND sg13g2_decap_8
XFILLER_28_260 VPWR VGND sg13g2_fill_2
XFILLER_28_282 VPWR VGND sg13g2_fill_2
XFILLER_43_263 VPWR VGND sg13g2_decap_8
XFILLER_16_499 VPWR VGND sg13g2_decap_4
XFILLER_32_937 VPWR VGND sg13g2_decap_8
XFILLER_32_948 VPWR VGND sg13g2_decap_8
XFILLER_40_970 VPWR VGND sg13g2_decap_8
XFILLER_7_120 VPWR VGND sg13g2_fill_2
XFILLER_11_193 VPWR VGND sg13g2_fill_1
X_3320_ _1050_ videogen.fancy_shader.video_y\[4\] videogen.fancy_shader.n646\[4\]
+ VPWR VGND sg13g2_nand2_1
X_3251_ net747 _0989_ _0362_ VPWR VGND sg13g2_nor2_1
XFILLER_26_1010 VPWR VGND sg13g2_decap_8
X_3182_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0914_ _0945_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_23_948 VPWR VGND sg13g2_decap_8
XFILLER_34_285 VPWR VGND sg13g2_decap_8
XFILLER_10_609 VPWR VGND sg13g2_decap_8
X_2966_ net608 net609 _0814_ VPWR VGND sg13g2_and2_1
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
X_4705_ _1994_ _1998_ _0613_ VPWR VGND sg13g2_nor2_1
X_2897_ _0784_ _0688_ _0717_ VPWR VGND sg13g2_nand2_2
X_4636_ net666 net717 _0189_ VPWR VGND sg13g2_nor2_1
X_5034__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_2_808 VPWR VGND sg13g2_fill_2
X_4567_ net681 net732 _0120_ VPWR VGND sg13g2_nor2_1
X_4498_ net652 net703 _0051_ VPWR VGND sg13g2_nor2_1
X_3518_ _1246_ _1247_ _1234_ _1248_ VPWR VGND sg13g2_nand3_1
X_5065__209 VPWR VGND net209 sg13g2_tiehi
X_3449_ _1178_ _1164_ _1165_ _1179_ VPWR VGND sg13g2_a21o_1
X_5119_ net799 VGND VPWR serialize.n427\[3\] serialize.n411\[1\] clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_27_78 VPWR VGND sg13g2_decap_8
XFILLER_14_915 VPWR VGND sg13g2_decap_8
XFILLER_13_425 VPWR VGND sg13g2_decap_4
XFILLER_40_244 VPWR VGND sg13g2_fill_2
XFILLER_22_970 VPWR VGND sg13g2_decap_8
XFILLER_5_679 VPWR VGND sg13g2_fill_2
XFILLER_4_156 VPWR VGND sg13g2_decap_4
XFILLER_4_38 VPWR VGND sg13g2_fill_1
XFILLER_49_834 VPWR VGND sg13g2_decap_8
XFILLER_48_311 VPWR VGND sg13g2_fill_1
XFILLER_1_874 VPWR VGND sg13g2_decap_8
XFILLER_48_344 VPWR VGND sg13g2_decap_8
X_2820_ _0703_ _0762_ _0767_ VPWR VGND sg13g2_nor2_2
XFILLER_9_952 VPWR VGND sg13g2_decap_8
X_2751_ _0750_ _0710_ _0713_ VPWR VGND sg13g2_nand2_2
X_2682_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\] net755 _0736_ _0553_
+ VPWR VGND sg13g2_mux2_1
X_4421_ _2111_ _2108_ _2109_ VPWR VGND sg13g2_xnor2_1
X_4352_ VGND VPWR _2019_ _2035_ _2047_ _2034_ sg13g2_a21oi_1
XFILLER_4_690 VPWR VGND sg13g2_fill_1
X_3303_ _1033_ _1027_ net546 VPWR VGND sg13g2_nand2_1
X_4283_ VGND VPWR _1985_ _1987_ _0505_ net570 sg13g2_a21oi_1
X_3234_ _0976_ _0977_ _0357_ VPWR VGND sg13g2_nor2_1
X_3165_ _0934_ net628 _0933_ VPWR VGND sg13g2_xnor2_1
X_3096_ _0878_ _0880_ _0883_ _0886_ VPWR VGND sg13g2_nor3_1
XFILLER_35_583 VPWR VGND sg13g2_decap_8
X_4860__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_23_734 VPWR VGND sg13g2_fill_2
X_3998_ _1619_ _1717_ _1722_ VPWR VGND sg13g2_and2_1
X_2949_ _0807_ _0802_ _0806_ _0801_ _0800_ VPWR VGND sg13g2_a22oi_1
X_4619_ net689 net741 _0172_ VPWR VGND sg13g2_nor2_1
XFILLER_49_119 VPWR VGND sg13g2_decap_4
XFILLER_16_1020 VPWR VGND sg13g2_decap_8
XFILLER_9_237 VPWR VGND sg13g2_fill_1
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_10_940 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_0_170 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_fill_1
X_4970_ net316 VGND VPWR _0517_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\]
+ _0165_ sg13g2_dfrbpq_1
X_3921_ _1640_ _1641_ _1646_ _1647_ VPWR VGND sg13g2_nor3_2
X_3852_ VGND VPWR _1581_ net2 videogen.test_lut_thingy.gol_counter_reg\[0\] sg13g2_or2_1
X_2803_ _0762_ _0679_ _0761_ VPWR VGND sg13g2_nand2_2
X_3783_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\] net582 _1513_ VPWR
+ VGND sg13g2_nor2_1
X_2734_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\] _0746_ _0511_
+ VPWR VGND sg13g2_mux2_1
X_4890__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_2665_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\] _0732_ _0566_
+ VPWR VGND sg13g2_mux2_1
X_2596_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\] _0704_ _0607_
+ VPWR VGND sg13g2_mux2_1
X_4404_ _2004_ _2093_ _2094_ _2095_ VPWR VGND sg13g2_nor3_1
X_4790__394 VPWR VGND net394 sg13g2_tiehi
X_4335_ _2031_ _2016_ _2029_ VPWR VGND sg13g2_nand2_1
XFILLER_5_92 VPWR VGND sg13g2_decap_4
X_4266_ _1962_ _1963_ _1969_ _1971_ _1972_ VPWR VGND sg13g2_nor4_1
X_3217_ net747 _0966_ _0351_ VPWR VGND sg13g2_nor2_1
XFILLER_28_804 VPWR VGND sg13g2_decap_4
X_4197_ VGND VPWR _0891_ _1913_ _1914_ _0647_ sg13g2_a21oi_1
XFILLER_39_185 VPWR VGND sg13g2_fill_1
X_3148_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0920_ _0922_ VPWR VGND
+ sg13g2_and2_1
X_3079_ _0869_ _0866_ _0868_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_870 VPWR VGND sg13g2_fill_1
XFILLER_42_339 VPWR VGND sg13g2_decap_4
XFILLER_23_597 VPWR VGND sg13g2_decap_8
XFILLER_3_925 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_decap_8
Xfanout750 net751 net750 VPWR VGND sg13g2_buf_8
Xfanout772 net773 net772 VPWR VGND sg13g2_buf_8
Xfanout783 net792 net783 VPWR VGND sg13g2_buf_8
XFILLER_19_815 VPWR VGND sg13g2_decap_8
Xfanout761 ui_in[7] net761 VPWR VGND sg13g2_buf_8
Xfanout794 rst_n net794 VPWR VGND sg13g2_buf_8
XFILLER_18_358 VPWR VGND sg13g2_decap_8
XFILLER_18_369 VPWR VGND sg13g2_fill_1
XFILLER_33_306 VPWR VGND sg13g2_decap_8
XFILLER_14_564 VPWR VGND sg13g2_decap_8
X_4120_ VPWR _1843_ _1842_ VGND sg13g2_inv_1
X_4051_ _1768_ _1773_ _1762_ _1774_ VPWR VGND sg13g2_nand3_1
X_3002_ VGND VPWR serialize.n431\[5\] net699 net412 sg13g2_or2_1
XFILLER_49_483 VPWR VGND sg13g2_decap_8
XFILLER_37_667 VPWR VGND sg13g2_decap_8
XFILLER_25_807 VPWR VGND sg13g2_fill_2
X_4953_ net395 VGND VPWR _0500_ green_tmds_par\[9\] net646 sg13g2_dfrbpq_1
X_3904_ _1630_ net546 _1626_ VPWR VGND sg13g2_nand2_1
X_4884_ net228 VGND VPWR _0435_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\]
+ _0092_ sg13g2_dfrbpq_1
XFILLER_20_501 VPWR VGND sg13g2_fill_1
XFILLER_33_884 VPWR VGND sg13g2_decap_8
XFILLER_33_895 VPWR VGND sg13g2_fill_1
X_3835_ VGND VPWR _1564_ net575 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\]
+ sg13g2_or2_1
X_3766_ net620 _1490_ _1495_ _1496_ VPWR VGND sg13g2_nor3_1
X_4859__280 VPWR VGND net280 sg13g2_tiehi
X_2717_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\] _0743_ _0525_
+ VPWR VGND sg13g2_mux2_1
X_3697_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\] net579 _1427_ VPWR
+ VGND sg13g2_nor2_1
X_2648_ _0692_ _0695_ _0709_ _0727_ VPWR VGND sg13g2_nor3_2
X_2579_ _0694_ net619 _0674_ VPWR VGND sg13g2_xnor2_1
X_4318_ _2015_ tmds_green.dc_balancing_reg\[1\] net601 VPWR VGND sg13g2_nand2b_1
X_4249_ _1955_ _0653_ _1954_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_807 VPWR VGND sg13g2_fill_1
XFILLER_43_626 VPWR VGND sg13g2_decap_4
XFILLER_43_604 VPWR VGND sg13g2_fill_1
XFILLER_43_659 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_4
XFILLER_24_862 VPWR VGND sg13g2_decap_8
XFILLER_30_309 VPWR VGND sg13g2_decap_8
XFILLER_23_372 VPWR VGND sg13g2_fill_2
X_5038__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_7_505 VPWR VGND sg13g2_fill_1
XFILLER_2_265 VPWR VGND sg13g2_decap_8
Xfanout591 _0675_ net591 VPWR VGND sg13g2_buf_8
Xfanout580 net581 net580 VPWR VGND sg13g2_buf_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
XFILLER_46_464 VPWR VGND sg13g2_fill_2
XFILLER_33_114 VPWR VGND sg13g2_fill_1
XFILLER_34_637 VPWR VGND sg13g2_decap_8
XFILLER_14_350 VPWR VGND sg13g2_fill_1
XFILLER_33_169 VPWR VGND sg13g2_decap_8
XFILLER_30_821 VPWR VGND sg13g2_fill_2
X_3620_ _1301_ _1349_ net2 _1350_ VPWR VGND sg13g2_nand3_1
X_3551_ _1277_ _1278_ _1279_ _1280_ _1281_ VPWR VGND sg13g2_nor4_1
XFILLER_6_593 VPWR VGND sg13g2_fill_2
X_3482_ _1209_ _1207_ net544 _1212_ VPWR VGND sg13g2_a21o_1
X_4103_ VGND VPWR _1826_ _1825_ _1824_ sg13g2_or2_1
XFILLER_29_409 VPWR VGND sg13g2_decap_8
X_5083_ net248 VGND VPWR _0630_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\]
+ _0260_ sg13g2_dfrbpq_1
X_4034_ VPWR VGND _1755_ _1752_ _1754_ _1741_ _1757_ _1745_ sg13g2_a221oi_1
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
XFILLER_24_136 VPWR VGND sg13g2_fill_1
X_4936_ net402 VGND VPWR _0000_ videogen.mem_read net634 sg13g2_dfrbpq_2
X_4867_ net265 VGND VPWR _0418_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\]
+ _0075_ sg13g2_dfrbpq_1
XFILLER_21_898 VPWR VGND sg13g2_decap_4
X_3818_ _1548_ _1499_ _1547_ videogen.test_lut_thingy.gol_counter_reg\[3\] _0650_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_21_36 VPWR VGND sg13g2_fill_2
X_4798_ net378 VGND VPWR _0349_ videogen.fancy_shader.n646\[3\] net636 sg13g2_dfrbpq_1
X_3749_ _1475_ _1476_ _1477_ _1478_ _1479_ VPWR VGND sg13g2_nor4_1
XFILLER_43_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_fill_1
XFILLER_0_758 VPWR VGND sg13g2_decap_8
XFILLER_29_932 VPWR VGND sg13g2_decap_8
XFILLER_28_431 VPWR VGND sg13g2_fill_2
XFILLER_28_453 VPWR VGND sg13g2_decap_8
XFILLER_46_99 VPWR VGND sg13g2_fill_1
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_28_497 VPWR VGND sg13g2_fill_1
X_5079__369 VPWR VGND net369 sg13g2_tiehi
XFILLER_12_821 VPWR VGND sg13g2_decap_8
XFILLER_24_681 VPWR VGND sg13g2_fill_2
XFILLER_7_324 VPWR VGND sg13g2_decap_8
XFILLER_11_386 VPWR VGND sg13g2_fill_1
XFILLER_3_530 VPWR VGND sg13g2_fill_2
XFILLER_3_541 VPWR VGND sg13g2_fill_1
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_3_574 VPWR VGND sg13g2_decap_8
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_47_795 VPWR VGND sg13g2_fill_2
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_412 VPWR VGND sg13g2_decap_8
X_2982_ _0820_ _0827_ net18 VPWR VGND sg13g2_nor2b_1
XFILLER_15_670 VPWR VGND sg13g2_decap_8
X_4721_ net142 VGND VPWR _0272_ green_tmds_par\[1\] net646 sg13g2_dfrbpq_1
XFILLER_30_640 VPWR VGND sg13g2_fill_2
X_4652_ net684 net735 _0205_ VPWR VGND sg13g2_nor2_1
X_3603_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\] net572 _1333_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_30_695 VPWR VGND sg13g2_decap_4
X_4583_ net677 net729 _0136_ VPWR VGND sg13g2_nor2_1
X_3534_ net616 _1258_ _1263_ _1264_ VPWR VGND sg13g2_nor3_1
XFILLER_6_390 VPWR VGND sg13g2_fill_2
X_3465_ VPWR _1195_ _1194_ VGND sg13g2_inv_1
X_3396_ _1112_ _1125_ _1087_ _1126_ VPWR VGND sg13g2_nand3_1
X_5066_ net201 VGND VPWR _0613_ blue_tmds_par\[3\] net646 sg13g2_dfrbpq_1
XFILLER_29_228 VPWR VGND sg13g2_decap_4
XFILLER_38_784 VPWR VGND sg13g2_decap_4
X_4017_ _1740_ _1739_ _1736_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_401 VPWR VGND sg13g2_decap_4
XFILLER_26_968 VPWR VGND sg13g2_decap_8
XFILLER_40_415 VPWR VGND sg13g2_decap_4
X_4778__46 VPWR VGND net46 sg13g2_tiehi
XFILLER_40_459 VPWR VGND sg13g2_fill_1
XFILLER_12_128 VPWR VGND sg13g2_decap_4
X_4919_ net158 VGND VPWR _0470_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\]
+ _0127_ sg13g2_dfrbpq_1
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_555 VPWR VGND sg13g2_decap_8
XFILLER_48_548 VPWR VGND sg13g2_decap_8
XFILLER_17_935 VPWR VGND sg13g2_decap_8
XFILLER_16_456 VPWR VGND sg13g2_fill_1
XFILLER_32_916 VPWR VGND sg13g2_decap_8
XFILLER_43_286 VPWR VGND sg13g2_fill_1
XFILLER_25_990 VPWR VGND sg13g2_decap_8
XFILLER_31_448 VPWR VGND sg13g2_decap_8
XFILLER_31_459 VPWR VGND sg13g2_decap_8
XFILLER_4_850 VPWR VGND sg13g2_decap_4
XFILLER_4_894 VPWR VGND sg13g2_decap_8
X_3250_ _0989_ videogen.fancy_shader.video_y\[6\] _0988_ VPWR VGND sg13g2_xnor2_1
X_3181_ VGND VPWR _0944_ _0919_ _0916_ sg13g2_or2_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_47_592 VPWR VGND sg13g2_decap_8
XFILLER_35_710 VPWR VGND sg13g2_decap_4
XFILLER_35_743 VPWR VGND sg13g2_decap_8
XFILLER_23_927 VPWR VGND sg13g2_decap_8
XFILLER_34_297 VPWR VGND sg13g2_decap_4
X_4704_ net665 net716 _0257_ VPWR VGND sg13g2_nor2_1
X_2965_ _0671_ _0683_ _0813_ VPWR VGND sg13g2_and2_1
X_2896_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\] net786 _0783_ _0313_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_481 VPWR VGND sg13g2_decap_8
X_4635_ net666 net717 _0188_ VPWR VGND sg13g2_nor2_1
X_4934__255 VPWR VGND net255 sg13g2_tiehi
X_4566_ net683 net732 _0119_ VPWR VGND sg13g2_nor2_1
X_3517_ _1247_ net547 _1187_ VPWR VGND sg13g2_xnor2_1
X_4497_ net651 net702 _0050_ VPWR VGND sg13g2_nor2_1
X_3448_ _1178_ _1160_ _1169_ VPWR VGND sg13g2_nand2_1
X_3379_ videogen.fancy_shader.video_x\[9\] videogen.fancy_shader.n646\[9\] _1109_
+ VPWR VGND sg13g2_xor2_1
XFILLER_40_1019 VPWR VGND sg13g2_decap_8
X_5118_ net799 VGND VPWR serialize.n427\[2\] serialize.n411\[0\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_45_507 VPWR VGND sg13g2_fill_1
XFILLER_38_592 VPWR VGND sg13g2_decap_8
X_5049_ net130 VGND VPWR _0596_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\]
+ _0244_ sg13g2_dfrbpq_1
XFILLER_25_231 VPWR VGND sg13g2_fill_2
XFILLER_5_636 VPWR VGND sg13g2_fill_1
XFILLER_5_658 VPWR VGND sg13g2_decap_8
XFILLER_1_853 VPWR VGND sg13g2_decap_8
XFILLER_49_824 VPWR VGND sg13g2_fill_1
XFILLER_48_323 VPWR VGND sg13g2_decap_8
XFILLER_0_374 VPWR VGND sg13g2_fill_1
XFILLER_0_396 VPWR VGND sg13g2_fill_2
XFILLER_44_573 VPWR VGND sg13g2_decap_4
XFILLER_16_297 VPWR VGND sg13g2_decap_8
XFILLER_32_779 VPWR VGND sg13g2_decap_8
XFILLER_9_931 VPWR VGND sg13g2_decap_8
XFILLER_12_470 VPWR VGND sg13g2_fill_1
XFILLER_13_993 VPWR VGND sg13g2_decap_8
X_2750_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\] net782 _0749_ _0489_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_289 VPWR VGND sg13g2_decap_8
X_4765__71 VPWR VGND net71 sg13g2_tiehi
X_2681_ _0723_ _0731_ _0736_ VPWR VGND sg13g2_nor2b_2
XFILLER_8_463 VPWR VGND sg13g2_fill_1
XFILLER_8_452 VPWR VGND sg13g2_decap_8
X_4420_ _2110_ _2109_ _2108_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_496 VPWR VGND sg13g2_decap_8
X_4351_ _2046_ _2043_ _2044_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_190 VPWR VGND sg13g2_decap_4
X_3302_ VGND VPWR _1032_ net546 _1027_ sg13g2_or2_1
X_4282_ VGND VPWR _0885_ _1982_ _1987_ _1986_ sg13g2_a21oi_1
X_3233_ net803 VPWR _0977_ VGND net608 _0974_ sg13g2_o21ai_1
X_3164_ _0931_ _0932_ _0933_ VPWR VGND sg13g2_nor2_1
X_3095_ _0884_ net548 _0885_ VPWR VGND sg13g2_nor2b_2
XFILLER_35_540 VPWR VGND sg13g2_fill_1
XFILLER_23_757 VPWR VGND sg13g2_decap_8
X_3997_ _1719_ _1721_ _1716_ _0376_ VPWR VGND sg13g2_nand3_1
X_2948_ _0806_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] _0804_ _0805_
+ VPWR VGND sg13g2_and3_1
X_2879_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\] net762 _0780_ _0391_
+ VPWR VGND sg13g2_mux2_1
X_4618_ net689 net741 _0171_ VPWR VGND sg13g2_nor2_1
X_4549_ net679 net730 _0102_ VPWR VGND sg13g2_nor2_1
XFILLER_45_337 VPWR VGND sg13g2_fill_2
X_5006__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_14_757 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_4
XFILLER_10_996 VPWR VGND sg13g2_decap_8
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_5_433 VPWR VGND sg13g2_fill_1
XFILLER_5_488 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_4
XFILLER_1_683 VPWR VGND sg13g2_decap_4
XFILLER_23_1025 VPWR VGND sg13g2_decap_4
X_3920_ _1637_ _1641_ _1643_ _1646_ VPWR VGND sg13g2_nor3_1
XFILLER_17_551 VPWR VGND sg13g2_decap_8
XFILLER_44_381 VPWR VGND sg13g2_decap_4
XFILLER_32_510 VPWR VGND sg13g2_decap_8
XFILLER_32_521 VPWR VGND sg13g2_decap_8
X_4994__219 VPWR VGND net219 sg13g2_tiehi
X_3851_ _1579_ VPWR _1580_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\]
+ net580 sg13g2_o21ai_1
XFILLER_32_576 VPWR VGND sg13g2_decap_8
X_3782_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\] net559 _1512_ VPWR
+ VGND sg13g2_nor2_1
X_2802_ _0673_ VPWR _0761_ VGND _0682_ _0684_ sg13g2_o21ai_1
X_2733_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\] _0746_ _0512_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_1007 VPWR VGND sg13g2_decap_8
XFILLER_8_282 VPWR VGND sg13g2_decap_8
XFILLER_8_260 VPWR VGND sg13g2_decap_8
X_2664_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\] _0732_ _0567_
+ VPWR VGND sg13g2_mux2_1
X_2595_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\] _0704_ _0608_
+ VPWR VGND sg13g2_mux2_1
X_4403_ _2094_ _2074_ _2091_ VPWR VGND sg13g2_xnor2_1
X_4334_ _2016_ _2029_ _2030_ VPWR VGND sg13g2_and2_1
X_4265_ _0890_ _1970_ _1971_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_131 VPWR VGND sg13g2_decap_8
X_3216_ _0966_ videogen.fancy_shader.n646\[5\] _0965_ VPWR VGND sg13g2_xnor2_1
X_4196_ _0860_ tmds_red.n114 _1913_ VPWR VGND sg13g2_xor2_1
X_3147_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0920_ _0921_ VPWR VGND
+ sg13g2_nor2_1
XFILLER_28_838 VPWR VGND sg13g2_decap_8
XFILLER_43_819 VPWR VGND sg13g2_decap_8
XFILLER_39_1021 VPWR VGND sg13g2_decap_8
X_3078_ VGND VPWR _0854_ net548 _0868_ _0867_ sg13g2_a21oi_1
XFILLER_11_716 VPWR VGND sg13g2_decap_4
XFILLER_23_576 VPWR VGND sg13g2_fill_1
XFILLER_7_709 VPWR VGND sg13g2_decap_8
XFILLER_40_13 VPWR VGND sg13g2_fill_2
XFILLER_3_904 VPWR VGND sg13g2_decap_8
XFILLER_2_414 VPWR VGND sg13g2_decap_4
XFILLER_49_77 VPWR VGND sg13g2_decap_8
Xfanout751 _0648_ net751 VPWR VGND sg13g2_buf_8
Xfanout740 net742 net740 VPWR VGND sg13g2_buf_8
Xfanout773 net776 net773 VPWR VGND sg13g2_buf_8
Xfanout762 net766 net762 VPWR VGND sg13g2_buf_8
Xfanout784 net786 net784 VPWR VGND sg13g2_buf_8
XFILLER_18_326 VPWR VGND sg13g2_decap_4
Xfanout795 net803 net795 VPWR VGND sg13g2_buf_8
XFILLER_14_532 VPWR VGND sg13g2_fill_2
XFILLER_26_392 VPWR VGND sg13g2_decap_4
XFILLER_14_587 VPWR VGND sg13g2_fill_2
XFILLER_41_395 VPWR VGND sg13g2_fill_1
XFILLER_10_760 VPWR VGND sg13g2_fill_1
XFILLER_5_230 VPWR VGND sg13g2_decap_8
XFILLER_49_440 VPWR VGND sg13g2_decap_4
X_4050_ _1773_ _1771_ _1772_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_462 VPWR VGND sg13g2_decap_8
X_3001_ net699 net412 serialize.n431\[4\] VPWR VGND sg13g2_nor2b_1
XFILLER_37_635 VPWR VGND sg13g2_fill_1
X_4952_ net397 VGND VPWR _0499_ green_tmds_par\[8\] net642 sg13g2_dfrbpq_1
X_4883_ net230 VGND VPWR _0434_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\]
+ _0091_ sg13g2_dfrbpq_1
X_3903_ _1627_ _1628_ _1629_ VPWR VGND sg13g2_and2_1
XFILLER_33_852 VPWR VGND sg13g2_decap_8
XFILLER_33_863 VPWR VGND sg13g2_fill_2
X_3834_ _1563_ _0674_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_32_373 VPWR VGND sg13g2_decap_8
X_3765_ _1491_ _1492_ _1493_ _1494_ _1495_ VPWR VGND sg13g2_nor4_1
X_3696_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\] net566 _1426_ VPWR
+ VGND sg13g2_nor2_1
X_2716_ _0743_ _0702_ _0706_ VPWR VGND sg13g2_nand2_2
X_2647_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\] net789 _0726_ _0578_
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_16 VPWR VGND sg13g2_decap_8
X_2578_ _0693_ net543 _0691_ VPWR VGND sg13g2_nand2_1
X_4317_ _0618_ net797 _2005_ _2014_ VPWR VGND sg13g2_and3_1
X_4248_ _0883_ VPWR _1954_ VGND _0878_ _0880_ sg13g2_o21ai_1
X_4179_ _1548_ _1620_ _1902_ VPWR VGND net1 sg13g2_nand3b_1
XFILLER_28_679 VPWR VGND sg13g2_decap_8
XFILLER_27_178 VPWR VGND sg13g2_decap_8
XFILLER_35_79 VPWR VGND sg13g2_fill_1
XFILLER_11_524 VPWR VGND sg13g2_decap_8
X_4838__321 VPWR VGND net321 sg13g2_tiehi
XFILLER_3_723 VPWR VGND sg13g2_decap_8
XFILLER_2_211 VPWR VGND sg13g2_fill_1
XFILLER_2_299 VPWR VGND sg13g2_fill_2
Xfanout570 net571 net570 VPWR VGND sg13g2_buf_8
Xfanout592 net595 net592 VPWR VGND sg13g2_buf_8
Xfanout581 _0690_ net581 VPWR VGND sg13g2_buf_8
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_46_443 VPWR VGND sg13g2_fill_1
XFILLER_46_432 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_668 VPWR VGND sg13g2_decap_8
XFILLER_30_888 VPWR VGND sg13g2_decap_8
X_3550_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\] net577 _1280_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_6_572 VPWR VGND sg13g2_decap_8
X_3481_ _1207_ VPWR _1211_ VGND _1206_ _1210_ sg13g2_o21ai_1
X_4102_ _1813_ _1818_ _1825_ VPWR VGND sg13g2_nor2_1
X_5082_ net283 VGND VPWR _0629_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\]
+ _0259_ sg13g2_dfrbpq_1
X_4033_ _1755_ _1754_ _1746_ _1756_ VPWR VGND sg13g2_a21o_1
XFILLER_25_605 VPWR VGND sg13g2_decap_4
XFILLER_25_649 VPWR VGND sg13g2_fill_2
X_4935_ net256 VGND VPWR _0003_ videogen.test_lut_thingy.pixel_feeder_inst.state\[1\]
+ net634 sg13g2_dfrbpq_1
XFILLER_21_800 VPWR VGND sg13g2_decap_4
X_4866_ net267 VGND VPWR _0417_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\]
+ _0074_ sg13g2_dfrbpq_1
X_4947__41 VPWR VGND net41 sg13g2_tiehi
X_4797_ net380 VGND VPWR _0348_ videogen.fancy_shader.n646\[2\] net637 sg13g2_dfrbpq_2
XFILLER_21_877 VPWR VGND sg13g2_decap_8
X_3817_ _0650_ _1546_ _1547_ VPWR VGND sg13g2_nor2_1
X_3748_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\] net582 _1478_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_21_59 VPWR VGND sg13g2_fill_2
X_3679_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\] net553 _1409_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_737 VPWR VGND sg13g2_decap_8
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_911 VPWR VGND sg13g2_decap_8
XFILLER_47_229 VPWR VGND sg13g2_fill_2
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_29_988 VPWR VGND sg13g2_decap_8
XFILLER_16_627 VPWR VGND sg13g2_fill_2
XFILLER_43_468 VPWR VGND sg13g2_decap_8
X_4805__364 VPWR VGND net364 sg13g2_tiehi
XFILLER_24_660 VPWR VGND sg13g2_decap_8
XFILLER_11_310 VPWR VGND sg13g2_decap_4
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_30_129 VPWR VGND sg13g2_fill_1
XFILLER_7_17 VPWR VGND sg13g2_decap_4
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_8_848 VPWR VGND sg13g2_decap_4
X_5049__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_46_251 VPWR VGND sg13g2_decap_4
XFILLER_19_443 VPWR VGND sg13g2_fill_1
XFILLER_34_457 VPWR VGND sg13g2_fill_2
XFILLER_43_991 VPWR VGND sg13g2_decap_8
X_2981_ _0818_ VPWR _0827_ VGND _0825_ _0826_ sg13g2_o21ai_1
XFILLER_22_619 VPWR VGND sg13g2_decap_8
XFILLER_42_490 VPWR VGND sg13g2_decap_8
X_4720_ net143 VGND VPWR _0271_ green_tmds_par\[0\] net646 sg13g2_dfrbpq_1
X_4651_ net669 net719 _0204_ VPWR VGND sg13g2_nor2_1
XFILLER_30_663 VPWR VGND sg13g2_fill_2
X_3602_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\] net559 _1332_ VPWR
+ VGND sg13g2_nor2_1
X_4582_ net677 net728 _0135_ VPWR VGND sg13g2_nor2_1
X_3533_ _1259_ _1260_ _1261_ _1262_ _1263_ VPWR VGND sg13g2_nor4_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_3464_ VGND VPWR _1194_ _1193_ _1192_ sg13g2_or2_1
X_3395_ _1125_ _1120_ _1124_ VPWR VGND sg13g2_nand2_1
X_5065_ net209 VGND VPWR _0612_ blue_tmds_par\[2\] net641 sg13g2_dfrbpq_1
X_4016_ _1739_ _1639_ _1738_ VPWR VGND sg13g2_xnor2_1
X_4828__331 VPWR VGND net331 sg13g2_tiehi
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_25_413 VPWR VGND sg13g2_decap_8
XFILLER_26_947 VPWR VGND sg13g2_decap_8
XFILLER_37_295 VPWR VGND sg13g2_decap_8
X_5019__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_13_619 VPWR VGND sg13g2_decap_8
X_4918_ net160 VGND VPWR _0469_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\]
+ _0126_ sg13g2_dfrbpq_1
XFILLER_21_652 VPWR VGND sg13g2_fill_1
X_4849_ net299 VGND VPWR _0400_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\]
+ _0057_ sg13g2_dfrbpq_1
XFILLER_21_696 VPWR VGND sg13g2_decap_8
XFILLER_5_829 VPWR VGND sg13g2_fill_1
X_4835__324 VPWR VGND net324 sg13g2_tiehi
X_4870__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_0_534 VPWR VGND sg13g2_decap_8
XFILLER_48_527 VPWR VGND sg13g2_decap_8
XFILLER_29_741 VPWR VGND sg13g2_fill_1
XFILLER_29_752 VPWR VGND sg13g2_fill_1
XFILLER_29_796 VPWR VGND sg13g2_decap_8
XFILLER_12_696 VPWR VGND sg13g2_decap_4
X_3180_ _0793_ _0943_ _0329_ VPWR VGND sg13g2_nor2_1
XFILLER_39_549 VPWR VGND sg13g2_fill_1
XFILLER_39_527 VPWR VGND sg13g2_decap_8
XFILLER_19_240 VPWR VGND sg13g2_fill_1
XFILLER_47_571 VPWR VGND sg13g2_decap_8
XFILLER_23_906 VPWR VGND sg13g2_decap_8
XFILLER_35_766 VPWR VGND sg13g2_decap_4
XFILLER_34_254 VPWR VGND sg13g2_fill_1
X_2964_ VGND VPWR _0649_ net15 _0684_ _0671_ sg13g2_a21oi_2
X_4703_ net662 net713 _0256_ VPWR VGND sg13g2_nor2_1
X_2895_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\] net776 _0783_ _0314_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_983 VPWR VGND sg13g2_decap_8
X_4634_ net670 net721 _0187_ VPWR VGND sg13g2_nor2_1
X_4565_ net681 net732 _0118_ VPWR VGND sg13g2_nor2_1
X_3516_ _1245_ VPWR _1246_ VGND _1242_ _1243_ sg13g2_o21ai_1
X_4496_ net651 net702 _0049_ VPWR VGND sg13g2_nor2_1
X_3447_ _1177_ _1174_ _1175_ VPWR VGND sg13g2_xnor2_1
X_3378_ _1100_ VPWR _1108_ VGND _1105_ _1106_ sg13g2_o21ai_1
X_5117_ net799 VGND VPWR serialize.n427\[1\] serialize.n452 clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5048_ net157 VGND VPWR _0595_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\]
+ _0243_ sg13g2_dfrbpq_1
XFILLER_26_766 VPWR VGND sg13g2_decap_8
XFILLER_26_777 VPWR VGND sg13g2_fill_2
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_40_213 VPWR VGND sg13g2_fill_2
XFILLER_25_287 VPWR VGND sg13g2_decap_8
XFILLER_43_68 VPWR VGND sg13g2_fill_2
X_4759__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_21_460 VPWR VGND sg13g2_fill_1
XFILLER_49_1023 VPWR VGND sg13g2_decap_4
XFILLER_1_832 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_4
XFILLER_49_869 VPWR VGND sg13g2_decap_8
XFILLER_36_508 VPWR VGND sg13g2_fill_2
XFILLER_48_379 VPWR VGND sg13g2_decap_8
XFILLER_1_1014 VPWR VGND sg13g2_decap_8
XFILLER_16_210 VPWR VGND sg13g2_decap_8
XFILLER_29_593 VPWR VGND sg13g2_decap_8
XFILLER_44_552 VPWR VGND sg13g2_decap_8
XFILLER_16_265 VPWR VGND sg13g2_decap_8
XFILLER_31_213 VPWR VGND sg13g2_decap_8
XFILLER_31_235 VPWR VGND sg13g2_decap_8
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_13_972 VPWR VGND sg13g2_decap_8
XFILLER_31_268 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_fill_1
XFILLER_12_482 VPWR VGND sg13g2_decap_8
XFILLER_31_279 VPWR VGND sg13g2_fill_2
XFILLER_9_987 VPWR VGND sg13g2_decap_8
XFILLER_12_493 VPWR VGND sg13g2_fill_1
X_5021__43 VPWR VGND net43 sg13g2_tiehi
X_2680_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\] _0735_ _0554_
+ VPWR VGND sg13g2_mux2_1
X_4818__341 VPWR VGND net341 sg13g2_tiehi
X_4780__42 VPWR VGND net42 sg13g2_tiehi
X_4350_ _2042_ _2044_ _2045_ VPWR VGND sg13g2_nor2_1
X_3301_ _1031_ _1029_ _1030_ VPWR VGND sg13g2_xnor2_1
X_4281_ _1918_ _1977_ _1986_ VPWR VGND sg13g2_nor2_1
X_3232_ net608 _0974_ _0976_ VPWR VGND sg13g2_and2_1
X_3163_ _0932_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] _0792_ VPWR
+ VGND sg13g2_nand2_1
X_3094_ _0884_ _0881_ _0883_ _0856_ _0652_ VPWR VGND sg13g2_a22oi_1
X_4825__334 VPWR VGND net334 sg13g2_tiehi
XFILLER_23_736 VPWR VGND sg13g2_fill_1
XFILLER_22_268 VPWR VGND sg13g2_fill_2
X_3996_ VGND VPWR _1721_ _1720_ _1718_ sg13g2_or2_1
X_2947_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ _0805_ VPWR VGND sg13g2_nor2_1
X_4617_ net689 net741 _0170_ VPWR VGND sg13g2_nor2_1
X_4756__83 VPWR VGND net83 sg13g2_tiehi
X_2878_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\] net752 _0780_ _0392_
+ VPWR VGND sg13g2_mux2_1
X_4548_ net655 net706 _0101_ VPWR VGND sg13g2_nor2_1
X_4832__327 VPWR VGND net327 sg13g2_tiehi
X_4479_ net662 net713 _0032_ VPWR VGND sg13g2_nor2_1
X_5069__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_38_35 VPWR VGND sg13g2_decap_8
X_4869__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_46_817 VPWR VGND sg13g2_decap_4
XFILLER_14_725 VPWR VGND sg13g2_fill_2
X_4876__243 VPWR VGND net243 sg13g2_tiehi
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_10_975 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_1_662 VPWR VGND sg13g2_decap_8
X_4848__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_23_1004 VPWR VGND sg13g2_decap_8
XFILLER_49_644 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_decap_4
XFILLER_36_327 VPWR VGND sg13g2_fill_1
XFILLER_45_894 VPWR VGND sg13g2_decap_8
X_3850_ _1576_ _1577_ _1578_ _1579_ VPWR VGND sg13g2_nor3_1
X_3781_ net614 VPWR _1511_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[3\]
+ net572 sg13g2_o21ai_1
X_2801_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\] _0760_ _0449_
+ VPWR VGND sg13g2_mux2_1
X_2732_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\] _0746_ _0513_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_740 VPWR VGND sg13g2_fill_1
XFILLER_9_795 VPWR VGND sg13g2_decap_4
XFILLER_8_294 VPWR VGND sg13g2_fill_2
X_2663_ net762 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\] _0732_ _0568_
+ VPWR VGND sg13g2_mux2_1
X_2594_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\] _0704_ _0609_
+ VPWR VGND sg13g2_mux2_1
X_4402_ net604 _2074_ _2093_ VPWR VGND sg13g2_nor2_1
X_4753__86 VPWR VGND net86 sg13g2_tiehi
X_4333_ _2027_ tmds_green.dc_balancing_reg\[2\] _2029_ VPWR VGND sg13g2_xor2_1
X_4264_ _1945_ _1965_ _1970_ VPWR VGND sg13g2_nor2_1
XFILLER_39_110 VPWR VGND sg13g2_decap_8
X_3215_ net751 _0964_ _0965_ _0350_ VPWR VGND sg13g2_nor3_1
X_4195_ VGND VPWR net607 _1912_ _0384_ net750 sg13g2_a21oi_1
XFILLER_39_165 VPWR VGND sg13g2_fill_1
X_3146_ _0917_ _0919_ _0920_ _0318_ VPWR VGND sg13g2_nor3_1
X_3077_ tmds_red.n126 tmds_red.n132 _0867_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_1000 VPWR VGND sg13g2_decap_8
XFILLER_23_500 VPWR VGND sg13g2_fill_1
XFILLER_36_894 VPWR VGND sg13g2_decap_4
XFILLER_23_555 VPWR VGND sg13g2_decap_8
XFILLER_11_728 VPWR VGND sg13g2_fill_2
X_3979_ VGND VPWR _1625_ _1701_ _1705_ _1704_ sg13g2_a21oi_1
XFILLER_46_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_56 VPWR VGND sg13g2_decap_8
Xfanout730 net731 net730 VPWR VGND sg13g2_buf_8
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
Xfanout774 net775 net774 VPWR VGND sg13g2_buf_8
Xfanout752 net753 net752 VPWR VGND sg13g2_buf_8
Xfanout785 net786 net785 VPWR VGND sg13g2_buf_1
Xfanout763 net766 net763 VPWR VGND sg13g2_buf_1
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_8
XFILLER_27_850 VPWR VGND sg13g2_decap_4
X_5075__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_14_500 VPWR VGND sg13g2_fill_2
XFILLER_26_360 VPWR VGND sg13g2_decap_4
XFILLER_6_721 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
X_4815__344 VPWR VGND net344 sg13g2_tiehi
XFILLER_2_993 VPWR VGND sg13g2_decap_8
X_3000_ net700 net411 serialize.n431\[3\] VPWR VGND sg13g2_nor2b_1
XFILLER_36_102 VPWR VGND sg13g2_fill_2
XFILLER_25_809 VPWR VGND sg13g2_fill_1
XFILLER_36_157 VPWR VGND sg13g2_decap_8
XFILLER_36_168 VPWR VGND sg13g2_fill_2
X_4951_ net399 VGND VPWR _0498_ green_tmds_par\[6\] net644 sg13g2_dfrbpq_1
XFILLER_18_883 VPWR VGND sg13g2_decap_8
X_4882_ net232 VGND VPWR _0433_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\]
+ _0090_ sg13g2_dfrbpq_1
XFILLER_17_393 VPWR VGND sg13g2_decap_4
X_3902_ VGND VPWR _1628_ _1626_ _1036_ sg13g2_or2_1
X_4822__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_20_514 VPWR VGND sg13g2_decap_8
X_3833_ VGND VPWR _1562_ net562 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\]
+ sg13g2_or2_1
X_3764_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\] net584 _1494_ VPWR
+ VGND sg13g2_nor2_1
X_3695_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\] net556 _1425_ VPWR
+ VGND sg13g2_nor2_1
X_2715_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\] _0742_ _0526_
+ VPWR VGND sg13g2_mux2_1
X_2646_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\] net775 _0726_ _0579_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_919 VPWR VGND sg13g2_decap_8
X_2577_ net543 _0691_ _0692_ VPWR VGND sg13g2_and2_1
X_4316_ _2013_ VPWR _2014_ VGND tmds_blue.vsync _1999_ sg13g2_o21ai_1
X_4247_ VGND VPWR _1930_ _1938_ _1953_ _1937_ sg13g2_a21oi_1
X_4178_ VGND VPWR _1901_ _1449_ _1352_ sg13g2_or2_1
X_3129_ _0898_ _0906_ _0907_ _0310_ VPWR VGND sg13g2_nor3_1
XFILLER_23_341 VPWR VGND sg13g2_decap_8
XFILLER_24_842 VPWR VGND sg13g2_decap_8
XFILLER_11_503 VPWR VGND sg13g2_decap_8
XFILLER_23_352 VPWR VGND sg13g2_fill_2
XFILLER_24_897 VPWR VGND sg13g2_decap_8
XFILLER_11_558 VPWR VGND sg13g2_decap_4
XFILLER_23_385 VPWR VGND sg13g2_fill_2
XFILLER_13_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_289 VPWR VGND sg13g2_decap_4
Xfanout560 net568 net560 VPWR VGND sg13g2_buf_1
Xfanout571 _0837_ net571 VPWR VGND sg13g2_buf_8
Xfanout582 net583 net582 VPWR VGND sg13g2_buf_8
Xfanout593 net595 net593 VPWR VGND sg13g2_buf_1
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_19_636 VPWR VGND sg13g2_decap_8
XFILLER_46_477 VPWR VGND sg13g2_decap_8
XFILLER_46_466 VPWR VGND sg13g2_fill_1
X_4728__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_15_842 VPWR VGND sg13g2_decap_8
XFILLER_15_886 VPWR VGND sg13g2_decap_8
XFILLER_25_91 VPWR VGND sg13g2_decap_4
XFILLER_30_845 VPWR VGND sg13g2_decap_8
X_3480_ net544 _1203_ _1209_ _1210_ VPWR VGND sg13g2_nor3_1
XFILLER_44_4 VPWR VGND sg13g2_fill_1
X_4101_ VPWR VGND _1811_ _1814_ _1820_ _1816_ _1824_ _1817_ sg13g2_a221oi_1
X_5081_ net314 VGND VPWR _0628_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\]
+ _0258_ sg13g2_dfrbpq_1
XFILLER_38_912 VPWR VGND sg13g2_decap_8
X_4032_ _1745_ VPWR _1755_ VGND _1739_ _1741_ sg13g2_o21ai_1
XFILLER_2_95 VPWR VGND sg13g2_decap_4
XFILLER_25_628 VPWR VGND sg13g2_decap_8
X_4934_ net255 VGND VPWR _0002_ videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ net635 sg13g2_dfrbpq_1
X_4865_ net268 VGND VPWR _0416_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\]
+ _0073_ sg13g2_dfrbpq_1
XFILLER_32_193 VPWR VGND sg13g2_fill_1
XFILLER_20_355 VPWR VGND sg13g2_fill_1
X_4796_ net382 VGND VPWR _0347_ videogen.fancy_shader.n646\[1\] net649 sg13g2_dfrbpq_2
X_3816_ _0636_ _1522_ _1545_ _1546_ VPWR VGND sg13g2_nor3_1
X_3747_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\] net549 _1477_ VPWR
+ VGND sg13g2_nor2_1
X_3678_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\] net564 _1408_ VPWR
+ VGND sg13g2_nor2_1
X_2629_ _0680_ _0687_ _0720_ VPWR VGND sg13g2_nor2_2
XFILLER_0_716 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_29_967 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_28_488 VPWR VGND sg13g2_decap_8
XFILLER_15_127 VPWR VGND sg13g2_fill_1
XFILLER_24_683 VPWR VGND sg13g2_fill_1
XFILLER_8_827 VPWR VGND sg13g2_decap_4
XFILLER_11_344 VPWR VGND sg13g2_decap_4
X_4990__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_3_532 VPWR VGND sg13g2_fill_1
XFILLER_11_71 VPWR VGND sg13g2_fill_2
XFILLER_46_230 VPWR VGND sg13g2_decap_8
XFILLER_47_797 VPWR VGND sg13g2_fill_1
XFILLER_46_274 VPWR VGND sg13g2_decap_4
XFILLER_34_425 VPWR VGND sg13g2_decap_4
XFILLER_43_970 VPWR VGND sg13g2_decap_8
X_2980_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0822_ _0826_
+ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] sg13g2_a21oi_1
XFILLER_14_160 VPWR VGND sg13g2_decap_8
XFILLER_30_620 VPWR VGND sg13g2_fill_2
XFILLER_14_193 VPWR VGND sg13g2_decap_8
X_4650_ net668 net719 _0203_ VPWR VGND sg13g2_nor2_1
XFILLER_30_642 VPWR VGND sg13g2_fill_1
X_3601_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\] net549 _1331_ VPWR
+ VGND sg13g2_nor2_1
X_4581_ net676 net728 _0134_ VPWR VGND sg13g2_nor2_1
X_3532_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\] net554 _1262_ VPWR
+ VGND sg13g2_nor2_1
X_3463_ _1087_ _1191_ _1193_ VPWR VGND sg13g2_and2_1
XFILLER_6_392 VPWR VGND sg13g2_fill_1
X_3394_ _1124_ _1122_ _1123_ VPWR VGND sg13g2_xnor2_1
X_5064_ net217 VGND VPWR _0611_ blue_tmds_par\[1\] net646 sg13g2_dfrbpq_1
X_4015_ _1738_ _1122_ _1737_ VPWR VGND sg13g2_nand2_1
XFILLER_26_926 VPWR VGND sg13g2_decap_8
XFILLER_16_27 VPWR VGND sg13g2_decap_4
XFILLER_25_447 VPWR VGND sg13g2_decap_4
XFILLER_21_631 VPWR VGND sg13g2_decap_8
X_4917_ net162 VGND VPWR _0468_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\]
+ _0125_ sg13g2_dfrbpq_1
X_4848_ net301 VGND VPWR _0399_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[2\]
+ _0056_ sg13g2_dfrbpq_1
XFILLER_32_59 VPWR VGND sg13g2_decap_8
X_4779_ net44 VGND VPWR _0330_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\]
+ net631 sg13g2_dfrbpq_1
XFILLER_10_1017 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_43_277 VPWR VGND sg13g2_decap_8
X_4725__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_43_299 VPWR VGND sg13g2_decap_8
XFILLER_12_631 VPWR VGND sg13g2_decap_8
XFILLER_31_428 VPWR VGND sg13g2_fill_1
XFILLER_11_141 VPWR VGND sg13g2_decap_4
XFILLER_40_984 VPWR VGND sg13g2_decap_8
XFILLER_8_657 VPWR VGND sg13g2_decap_8
XFILLER_7_156 VPWR VGND sg13g2_decap_8
XFILLER_7_178 VPWR VGND sg13g2_fill_2
XFILLER_22_92 VPWR VGND sg13g2_decap_4
XFILLER_3_384 VPWR VGND sg13g2_decap_8
XFILLER_3_373 VPWR VGND sg13g2_fill_1
XFILLER_26_1024 VPWR VGND sg13g2_decap_4
XFILLER_19_263 VPWR VGND sg13g2_fill_1
X_4997__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_22_417 VPWR VGND sg13g2_decap_4
XFILLER_16_992 VPWR VGND sg13g2_decap_8
X_2963_ VGND VPWR _0649_ net14 _0682_ _0671_ sg13g2_a21oi_2
X_4702_ net665 net716 _0255_ VPWR VGND sg13g2_nor2_1
XFILLER_31_962 VPWR VGND sg13g2_decap_8
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
X_2894_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\] net766 _0783_ _0315_
+ VPWR VGND sg13g2_mux2_1
X_4633_ net670 net721 _0186_ VPWR VGND sg13g2_nor2_1
XFILLER_8_83 VPWR VGND sg13g2_fill_1
X_4564_ net681 net732 _0117_ VPWR VGND sg13g2_nor2_1
X_3515_ _1183_ _1244_ _1245_ VPWR VGND sg13g2_nor2b_1
X_4940__70 VPWR VGND net70 sg13g2_tiehi
X_4495_ net652 net703 _0048_ VPWR VGND sg13g2_nor2_1
X_3446_ _1175_ _1174_ _1176_ VPWR VGND sg13g2_xor2_1
X_3377_ videogen.fancy_shader.video_x\[8\] net610 _1107_ VPWR VGND sg13g2_xor2_1
X_5116_ net799 VGND VPWR serialize.n427\[0\] serialize.n450 clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5047_ net165 VGND VPWR _0594_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\]
+ _0242_ sg13g2_dfrbpq_1
XFILLER_27_26 VPWR VGND sg13g2_fill_1
XFILLER_27_48 VPWR VGND sg13g2_fill_2
XFILLER_25_211 VPWR VGND sg13g2_decap_8
XFILLER_26_756 VPWR VGND sg13g2_decap_4
X_4980__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_14_929 VPWR VGND sg13g2_decap_8
XFILLER_25_266 VPWR VGND sg13g2_fill_2
XFILLER_22_984 VPWR VGND sg13g2_decap_8
XFILLER_49_1002 VPWR VGND sg13g2_decap_8
XFILLER_1_811 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_fill_2
XFILLER_1_888 VPWR VGND sg13g2_decap_8
XFILLER_49_848 VPWR VGND sg13g2_decap_8
XFILLER_0_398 VPWR VGND sg13g2_fill_1
XFILLER_48_358 VPWR VGND sg13g2_decap_8
XFILLER_17_701 VPWR VGND sg13g2_fill_2
XFILLER_17_723 VPWR VGND sg13g2_decap_8
XFILLER_29_572 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_decap_4
XFILLER_16_233 VPWR VGND sg13g2_fill_2
XFILLER_17_767 VPWR VGND sg13g2_fill_2
XFILLER_17_789 VPWR VGND sg13g2_decap_8
XFILLER_32_715 VPWR VGND sg13g2_decap_8
XFILLER_32_737 VPWR VGND sg13g2_fill_1
XFILLER_13_951 VPWR VGND sg13g2_decap_8
XFILLER_12_461 VPWR VGND sg13g2_fill_1
XFILLER_8_443 VPWR VGND sg13g2_decap_4
XFILLER_9_966 VPWR VGND sg13g2_decap_8
X_3300_ VGND VPWR _1007_ _1009_ _1030_ _1008_ sg13g2_a21oi_1
XFILLER_4_682 VPWR VGND sg13g2_decap_4
XFILLER_3_170 VPWR VGND sg13g2_fill_1
X_4280_ _0884_ VPWR _1985_ VGND _1978_ _1984_ sg13g2_o21ai_1
X_5029__310 VPWR VGND net310 sg13g2_tiehi
X_3231_ _0974_ _0975_ _0356_ VPWR VGND sg13g2_nor2_1
X_3162_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0931_ VPWR VGND sg13g2_nor3_1
XFILLER_48_881 VPWR VGND sg13g2_decap_8
X_3093_ _0859_ _0882_ _0883_ VPWR VGND sg13g2_nor2_2
X_3995_ VGND VPWR _1720_ _1616_ _1449_ sg13g2_or2_1
X_2946_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\]
+ _0803_ _0804_ VPWR VGND sg13g2_nor3_2
X_2877_ _0728_ _0772_ _0780_ VPWR VGND sg13g2_nor2_2
X_4616_ net690 net744 _0169_ VPWR VGND sg13g2_nor2_1
X_4547_ net668 net720 _0100_ VPWR VGND sg13g2_nor2_1
X_4478_ net665 net716 _0031_ VPWR VGND sg13g2_nor2_1
X_3429_ net545 _1147_ _1159_ VPWR VGND sg13g2_nor2_1
XFILLER_39_870 VPWR VGND sg13g2_fill_1
XFILLER_26_575 VPWR VGND sg13g2_decap_8
XFILLER_41_567 VPWR VGND sg13g2_decap_4
XFILLER_10_954 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_fill_1
XFILLER_48_144 VPWR VGND sg13g2_decap_8
XFILLER_0_184 VPWR VGND sg13g2_decap_8
XFILLER_44_372 VPWR VGND sg13g2_decap_4
XFILLER_17_597 VPWR VGND sg13g2_decap_4
X_3780_ net621 _1504_ _1509_ _1510_ VPWR VGND sg13g2_nor3_1
X_2800_ net778 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\] _0760_ _0450_
+ VPWR VGND sg13g2_mux2_1
X_2731_ _0746_ _0706_ _0727_ VPWR VGND sg13g2_nand2_2
X_4738__115 VPWR VGND net115 sg13g2_tiehi
X_4401_ _2092_ _2074_ _2091_ VPWR VGND sg13g2_nand2b_1
X_2662_ net756 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\] _0732_ _0569_
+ VPWR VGND sg13g2_mux2_1
X_2593_ _0704_ _0688_ _0702_ VPWR VGND sg13g2_nand2_2
X_4332_ _2028_ _2027_ tmds_green.dc_balancing_reg\[2\] VPWR VGND sg13g2_nand2b_1
X_4263_ _0891_ _1946_ _1967_ _1968_ _1969_ VPWR VGND sg13g2_nor4_1
X_3214_ _0965_ videogen.fancy_shader.n646\[4\] net611 _0961_ VPWR VGND sg13g2_and3_2
X_4194_ _1912_ tmds_red.n102 _0891_ VPWR VGND sg13g2_xnor2_1
X_3145_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0916_ _0920_ VPWR VGND
+ sg13g2_and2_1
XFILLER_27_317 VPWR VGND sg13g2_fill_2
XFILLER_39_199 VPWR VGND sg13g2_fill_2
X_3076_ VGND VPWR _0857_ _0860_ _0866_ _0858_ sg13g2_a21oi_1
XFILLER_23_534 VPWR VGND sg13g2_fill_2
XFILLER_24_38 VPWR VGND sg13g2_decap_8
XFILLER_24_49 VPWR VGND sg13g2_fill_1
X_3978_ _1704_ _1699_ _1703_ VPWR VGND sg13g2_xnor2_1
X_2929_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\] _0790_ _0269_
+ VPWR VGND sg13g2_mux2_1
XFILLER_40_26 VPWR VGND sg13g2_decap_4
XFILLER_46_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_939 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
Xfanout731 net734 net731 VPWR VGND sg13g2_buf_2
Xfanout720 net724 net720 VPWR VGND sg13g2_buf_8
X_4986__250 VPWR VGND net250 sg13g2_tiehi
Xfanout742 net745 net742 VPWR VGND sg13g2_buf_8
Xfanout775 net776 net775 VPWR VGND sg13g2_buf_8
Xfanout753 net761 net753 VPWR VGND sg13g2_buf_8
Xfanout764 net765 net764 VPWR VGND sg13g2_buf_8
Xfanout797 net803 net797 VPWR VGND sg13g2_buf_8
Xfanout786 net792 net786 VPWR VGND sg13g2_buf_8
XFILLER_46_659 VPWR VGND sg13g2_fill_1
XFILLER_27_884 VPWR VGND sg13g2_decap_8
XFILLER_14_534 VPWR VGND sg13g2_fill_1
XFILLER_14_578 VPWR VGND sg13g2_fill_1
XFILLER_41_386 VPWR VGND sg13g2_decap_8
X_4958__385 VPWR VGND net385 sg13g2_tiehi
XFILLER_10_784 VPWR VGND sg13g2_decap_8
XFILLER_6_799 VPWR VGND sg13g2_fill_1
XFILLER_39_7 VPWR VGND sg13g2_decap_4
XFILLER_7_1010 VPWR VGND sg13g2_decap_8
XFILLER_2_972 VPWR VGND sg13g2_decap_8
XFILLER_1_460 VPWR VGND sg13g2_decap_4
XFILLER_37_604 VPWR VGND sg13g2_fill_2
XFILLER_49_497 VPWR VGND sg13g2_decap_8
X_5026__357 VPWR VGND net357 sg13g2_tiehi
X_4950_ net401 VGND VPWR _0497_ green_tmds_par\[2\] net644 sg13g2_dfrbpq_1
X_4881_ net233 VGND VPWR _0432_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\]
+ _0089_ sg13g2_dfrbpq_1
X_3901_ _1627_ _1036_ _1626_ VPWR VGND sg13g2_nand2_1
XFILLER_32_331 VPWR VGND sg13g2_fill_1
X_3832_ _1557_ _1558_ _1559_ _1560_ _1561_ VPWR VGND sg13g2_nor4_1
XFILLER_32_353 VPWR VGND sg13g2_fill_2
X_3763_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\] net562 _1493_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_560 VPWR VGND sg13g2_decap_8
XFILLER_20_559 VPWR VGND sg13g2_decap_8
X_3694_ net597 VPWR _1424_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\]
+ net590 sg13g2_o21ai_1
X_2714_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\] _0742_ _0527_
+ VPWR VGND sg13g2_mux2_1
X_2645_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\] net770 _0726_ _0580_
+ VPWR VGND sg13g2_mux2_1
X_2576_ net582 net572 _0691_ VPWR VGND sg13g2_and2_1
X_4315_ tmds_blue.vsync VPWR _2013_ VGND net606 hsync sg13g2_o21ai_1
X_4246_ net570 _1952_ _0503_ VPWR VGND sg13g2_nor2_1
X_4177_ _1894_ _1899_ _1795_ _1900_ VPWR VGND sg13g2_nand3_1
XFILLER_28_604 VPWR VGND sg13g2_fill_2
X_3128_ net629 _0800_ _0907_ VPWR VGND sg13g2_nor2_1
XFILLER_27_136 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_fill_2
X_3059_ net569 _0849_ _0273_ VPWR VGND sg13g2_nor2_1
XFILLER_24_821 VPWR VGND sg13g2_decap_8
XFILLER_35_180 VPWR VGND sg13g2_decap_4
XFILLER_24_876 VPWR VGND sg13g2_decap_8
XFILLER_2_246 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_decap_4
Xfanout550 net558 net550 VPWR VGND sg13g2_buf_1
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_19_615 VPWR VGND sg13g2_fill_1
Xfanout583 net591 net583 VPWR VGND sg13g2_buf_8
Xfanout572 net576 net572 VPWR VGND sg13g2_buf_8
Xfanout561 net562 net561 VPWR VGND sg13g2_buf_8
XFILLER_18_125 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
Xfanout594 net595 net594 VPWR VGND sg13g2_buf_8
XFILLER_46_456 VPWR VGND sg13g2_decap_4
XFILLER_14_342 VPWR VGND sg13g2_fill_2
XFILLER_25_70 VPWR VGND sg13g2_decap_4
X_5080_ net353 VGND VPWR _0627_ tmds_blue.dc_balancing_reg\[4\] net643 sg13g2_dfrbpq_2
X_4100_ _1822_ _1811_ _1823_ VPWR VGND sg13g2_nor2b_1
X_4031_ _1754_ _1740_ _1741_ VPWR VGND sg13g2_nand2_1
XFILLER_1_290 VPWR VGND sg13g2_fill_1
XFILLER_49_283 VPWR VGND sg13g2_fill_2
XFILLER_49_272 VPWR VGND sg13g2_decap_8
XFILLER_38_957 VPWR VGND sg13g2_fill_2
XFILLER_37_412 VPWR VGND sg13g2_decap_4
XFILLER_2_63 VPWR VGND sg13g2_decap_4
XFILLER_38_979 VPWR VGND sg13g2_decap_8
XFILLER_37_489 VPWR VGND sg13g2_decap_4
XFILLER_18_670 VPWR VGND sg13g2_fill_2
XFILLER_17_180 VPWR VGND sg13g2_decap_8
X_4933_ net254 VGND VPWR _0484_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\]
+ _0141_ sg13g2_dfrbpq_1
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
XFILLER_21_813 VPWR VGND sg13g2_decap_8
X_4864_ net270 VGND VPWR _0415_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\]
+ _0072_ sg13g2_dfrbpq_1
XFILLER_20_323 VPWR VGND sg13g2_fill_2
XFILLER_21_835 VPWR VGND sg13g2_decap_8
X_4902__192 VPWR VGND net192 sg13g2_tiehi
X_4795_ net384 VGND VPWR _0346_ videogen.fancy_shader.n646\[0\] net649 sg13g2_dfrbpq_2
X_3815_ net613 _1533_ _1544_ _1545_ VPWR VGND sg13g2_nor3_1
X_3746_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\] net559 _1476_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_367 VPWR VGND sg13g2_decap_4
X_4976__293 VPWR VGND net293 sg13g2_tiehi
X_3677_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\] net577 _1407_ VPWR
+ VGND sg13g2_nor2_1
X_2628_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\] _0719_ _0590_
+ VPWR VGND sg13g2_mux2_1
X_2559_ net625 net626 _0674_ VPWR VGND sg13g2_nor2_2
XFILLER_43_1019 VPWR VGND sg13g2_decap_8
X_4229_ VGND VPWR _0859_ _0875_ _1936_ _1934_ sg13g2_a21oi_1
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_946 VPWR VGND sg13g2_decap_8
XFILLER_16_629 VPWR VGND sg13g2_fill_1
XFILLER_37_990 VPWR VGND sg13g2_decap_8
XFILLER_7_305 VPWR VGND sg13g2_decap_8
XFILLER_20_890 VPWR VGND sg13g2_decap_8
XFILLER_3_588 VPWR VGND sg13g2_decap_8
XFILLER_4_1013 VPWR VGND sg13g2_decap_8
XFILLER_34_459 VPWR VGND sg13g2_fill_1
XFILLER_42_481 VPWR VGND sg13g2_decap_4
XFILLER_15_684 VPWR VGND sg13g2_decap_4
X_4580_ net666 net717 _0133_ VPWR VGND sg13g2_nor2_1
X_3600_ net619 VPWR _1330_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\]
+ net582 sg13g2_o21ai_1
X_3531_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\] net563 _1261_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_7_883 VPWR VGND sg13g2_fill_2
X_4856__286 VPWR VGND net286 sg13g2_tiehi
X_3462_ VGND VPWR _1190_ _1191_ _1192_ _1087_ sg13g2_a21oi_1
X_3393_ _1123_ _1094_ _1096_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_0 VPWR VGND sg13g2_fill_2
X_5063_ net225 VGND VPWR _0610_ blue_tmds_par\[0\] net641 sg13g2_dfrbpq_1
XFILLER_38_721 VPWR VGND sg13g2_fill_2
XFILLER_38_765 VPWR VGND sg13g2_decap_4
XFILLER_38_754 VPWR VGND sg13g2_decap_8
X_4014_ _1103_ _1729_ _1737_ VPWR VGND sg13g2_and2_1
XFILLER_26_905 VPWR VGND sg13g2_decap_8
XFILLER_38_798 VPWR VGND sg13g2_decap_8
XFILLER_16_39 VPWR VGND sg13g2_fill_2
XFILLER_41_919 VPWR VGND sg13g2_decap_8
X_4916_ net164 VGND VPWR _0467_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\]
+ _0124_ sg13g2_dfrbpq_1
XFILLER_34_993 VPWR VGND sg13g2_decap_8
X_4847_ net303 VGND VPWR _0398_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[1\]
+ _0055_ sg13g2_dfrbpq_1
XFILLER_32_38 VPWR VGND sg13g2_fill_2
XFILLER_33_492 VPWR VGND sg13g2_decap_4
XFILLER_20_153 VPWR VGND sg13g2_decap_8
X_4778_ net46 VGND VPWR _0329_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\]
+ net632 sg13g2_dfrbpq_2
XFILLER_20_186 VPWR VGND sg13g2_fill_2
X_3729_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\] net565 _1459_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_525 VPWR VGND sg13g2_decap_4
XFILLER_48_507 VPWR VGND sg13g2_fill_2
XFILLER_0_569 VPWR VGND sg13g2_decap_8
XFILLER_29_765 VPWR VGND sg13g2_decap_8
XFILLER_16_404 VPWR VGND sg13g2_decap_8
XFILLER_28_253 VPWR VGND sg13g2_decap_8
XFILLER_29_776 VPWR VGND sg13g2_fill_1
XFILLER_44_746 VPWR VGND sg13g2_fill_2
XFILLER_16_448 VPWR VGND sg13g2_fill_2
XFILLER_17_949 VPWR VGND sg13g2_decap_8
XFILLER_43_256 VPWR VGND sg13g2_decap_8
XFILLER_24_470 VPWR VGND sg13g2_fill_1
XFILLER_40_941 VPWR VGND sg13g2_fill_1
XFILLER_11_120 VPWR VGND sg13g2_decap_8
XFILLER_7_113 VPWR VGND sg13g2_decap_8
XFILLER_22_71 VPWR VGND sg13g2_decap_8
XFILLER_26_1003 VPWR VGND sg13g2_decap_8
X_4886__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_19_253 VPWR VGND sg13g2_decap_4
XFILLER_35_757 VPWR VGND sg13g2_fill_1
XFILLER_16_971 VPWR VGND sg13g2_decap_8
X_2962_ VGND VPWR _0649_ net13 _0678_ _0671_ sg13g2_a21oi_2
XFILLER_34_278 VPWR VGND sg13g2_decap_8
X_4701_ net661 net712 _0254_ VPWR VGND sg13g2_nor2_1
XFILLER_31_941 VPWR VGND sg13g2_decap_8
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
X_2893_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\] net755 _0783_ _0316_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_473 VPWR VGND sg13g2_decap_4
X_4632_ net688 net740 _0185_ VPWR VGND sg13g2_nor2_1
XFILLER_8_73 VPWR VGND sg13g2_fill_2
X_4563_ net682 net733 _0116_ VPWR VGND sg13g2_nor2_1
X_4494_ net651 net702 _0047_ VPWR VGND sg13g2_nor2_1
X_3514_ VGND VPWR _1244_ _1182_ _1179_ sg13g2_or2_1
X_3445_ _1013_ _1012_ _1175_ VPWR VGND sg13g2_xor2_1
X_3376_ net610 videogen.fancy_shader.video_x\[8\] _1106_ VPWR VGND sg13g2_nor2_1
X_5115_ net796 VGND VPWR _0262_ _0004_ clknet_3_2__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_38_540 VPWR VGND sg13g2_fill_1
X_5046_ net173 VGND VPWR _0593_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\]
+ _0241_ sg13g2_dfrbpq_1
X_5041__213 VPWR VGND net213 sg13g2_tiehi
XFILLER_40_215 VPWR VGND sg13g2_fill_1
XFILLER_40_204 VPWR VGND sg13g2_fill_1
XFILLER_40_259 VPWR VGND sg13g2_decap_4
XFILLER_22_963 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_fill_2
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_1_867 VPWR VGND sg13g2_decap_8
XFILLER_48_337 VPWR VGND sg13g2_decap_8
XFILLER_44_521 VPWR VGND sg13g2_decap_8
XFILLER_17_71 VPWR VGND sg13g2_decap_8
XFILLER_13_930 VPWR VGND sg13g2_decap_8
XFILLER_31_259 VPWR VGND sg13g2_fill_1
XFILLER_8_422 VPWR VGND sg13g2_decap_8
XFILLER_9_945 VPWR VGND sg13g2_decap_8
X_3230_ net795 VPWR _0975_ VGND net609 _0897_ sg13g2_o21ai_1
X_3161_ VPWR _0323_ _0930_ VGND sg13g2_inv_1
X_3092_ _0882_ _0865_ _0875_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_521 VPWR VGND sg13g2_fill_1
XFILLER_35_554 VPWR VGND sg13g2_decap_4
XFILLER_23_727 VPWR VGND sg13g2_decap_8
X_3994_ _0377_ _1716_ _1719_ VPWR VGND sg13g2_nand2_1
X_2945_ _0803_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\]
+ VPWR VGND sg13g2_nand2_1
X_2876_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\] net782 _0779_ _0393_
+ VPWR VGND sg13g2_mux2_1
X_4615_ net690 net743 _0168_ VPWR VGND sg13g2_nor2_1
X_4546_ net655 net706 _0099_ VPWR VGND sg13g2_nor2_1
X_4477_ net661 net712 _0030_ VPWR VGND sg13g2_nor2_1
X_3428_ _1158_ _1157_ _1156_ VPWR VGND sg13g2_nand2b_1
X_3359_ _1089_ videogen.fancy_shader.video_y\[8\] net610 VPWR VGND sg13g2_nand2_1
X_5029_ net310 VGND VPWR _0576_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\]
+ _0224_ sg13g2_dfrbpq_1
XFILLER_38_370 VPWR VGND sg13g2_decap_8
XFILLER_26_510 VPWR VGND sg13g2_decap_8
XFILLER_13_215 VPWR VGND sg13g2_fill_2
XFILLER_16_1013 VPWR VGND sg13g2_decap_8
XFILLER_10_933 VPWR VGND sg13g2_decap_8
XFILLER_21_270 VPWR VGND sg13g2_decap_4
XFILLER_22_782 VPWR VGND sg13g2_decap_8
X_4762__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_48_101 VPWR VGND sg13g2_decap_8
XFILLER_0_163 VPWR VGND sg13g2_decap_8
XFILLER_48_178 VPWR VGND sg13g2_fill_1
XFILLER_17_521 VPWR VGND sg13g2_decap_8
XFILLER_44_340 VPWR VGND sg13g2_decap_8
XFILLER_17_565 VPWR VGND sg13g2_decap_8
XFILLER_32_535 VPWR VGND sg13g2_decap_4
X_2730_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\] net790 _0745_ _0514_
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_292 VPWR VGND sg13g2_decap_8
X_2661_ _0732_ _0710_ _0731_ VPWR VGND sg13g2_nand2_2
XFILLER_8_296 VPWR VGND sg13g2_fill_1
XFILLER_8_274 VPWR VGND sg13g2_decap_4
X_4400_ _2089_ _2082_ _2091_ VPWR VGND sg13g2_xor2_1
X_2592_ _0674_ _0695_ videogen.mem_read _0703_ VPWR VGND sg13g2_nand3_1
XFILLER_5_981 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_fill_2
X_4331_ _2027_ _2024_ VPWR VGND _2022_ sg13g2_nand2b_2
XFILLER_5_96 VPWR VGND sg13g2_fill_1
XFILLER_5_85 VPWR VGND sg13g2_fill_2
X_4262_ _1965_ _1966_ _1968_ VPWR VGND sg13g2_nor2_1
X_3213_ VGND VPWR net611 _0961_ _0964_ videogen.fancy_shader.n646\[4\] sg13g2_a21oi_1
X_4193_ _1911_ net795 _1906_ _0383_ VPWR VGND sg13g2_a21o_1
X_3144_ _0919_ net793 _0918_ VPWR VGND sg13g2_nand2_2
XFILLER_28_808 VPWR VGND sg13g2_fill_2
XFILLER_48_690 VPWR VGND sg13g2_fill_2
X_3075_ _0865_ tmds_red.n100 _0859_ VPWR VGND sg13g2_nand2b_1
X_3977_ _1703_ _1675_ _1684_ VPWR VGND sg13g2_xnor2_1
X_4721__142 VPWR VGND net142 sg13g2_tiehi
X_2928_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\] _0790_ _0270_
+ VPWR VGND sg13g2_mux2_1
X_2859_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\] net768 _0776_ _0407_
+ VPWR VGND sg13g2_mux2_1
XFILLER_3_918 VPWR VGND sg13g2_decap_8
X_4529_ net658 net709 _0082_ VPWR VGND sg13g2_nor2_1
XFILLER_2_428 VPWR VGND sg13g2_fill_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
Xfanout721 net723 net721 VPWR VGND sg13g2_buf_8
Xfanout732 net733 net732 VPWR VGND sg13g2_buf_8
Xfanout710 net711 net710 VPWR VGND sg13g2_buf_8
X_4912__172 VPWR VGND net172 sg13g2_tiehi
Xfanout754 net755 net754 VPWR VGND sg13g2_buf_8
Xfanout743 net745 net743 VPWR VGND sg13g2_buf_8
Xfanout776 ui_in[5] net776 VPWR VGND sg13g2_buf_8
Xfanout765 net766 net765 VPWR VGND sg13g2_buf_8
Xfanout798 net802 net798 VPWR VGND sg13g2_buf_8
Xfanout787 net791 net787 VPWR VGND sg13g2_buf_8
XFILLER_42_822 VPWR VGND sg13g2_fill_1
XFILLER_14_546 VPWR VGND sg13g2_fill_1
XFILLER_26_384 VPWR VGND sg13g2_fill_2
XFILLER_6_756 VPWR VGND sg13g2_fill_1
XFILLER_2_951 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_36_104 VPWR VGND sg13g2_fill_1
X_4880_ net235 VGND VPWR _0431_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\]
+ _0088_ sg13g2_dfrbpq_1
X_3900_ _1010_ _1623_ _1626_ VPWR VGND sg13g2_nor2_2
X_3831_ net595 VPWR _1560_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\]
+ net579 sg13g2_o21ai_1
X_3762_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\] net574 _1492_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_387 VPWR VGND sg13g2_fill_2
X_2713_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\] _0742_ _0528_
+ VPWR VGND sg13g2_mux2_1
X_3693_ _0637_ _1411_ _1422_ _1423_ VPWR VGND sg13g2_nor3_1
X_2644_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\] net755 _0726_ _0581_
+ VPWR VGND sg13g2_mux2_1
X_2575_ _0690_ net624 net626 VPWR VGND sg13g2_nand2_2
X_4314_ VGND VPWR net605 net607 _0617_ _2000_ sg13g2_a21oi_1
XFILLER_19_17 VPWR VGND sg13g2_fill_2
X_4245_ VPWR VGND _1951_ _1949_ _1940_ _1919_ _1952_ _1939_ sg13g2_a221oi_1
X_4176_ _1898_ _1789_ _1792_ _1899_ VPWR VGND sg13g2_a21o_1
X_3127_ net629 _0800_ _0906_ VPWR VGND sg13g2_and2_1
XFILLER_43_619 VPWR VGND sg13g2_decap_8
XFILLER_42_118 VPWR VGND sg13g2_fill_2
XFILLER_35_27 VPWR VGND sg13g2_fill_2
X_3058_ _0849_ _0845_ _0848_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_387 VPWR VGND sg13g2_fill_1
XFILLER_2_258 VPWR VGND sg13g2_decap_8
Xfanout551 net552 net551 VPWR VGND sg13g2_buf_8
Xfanout573 net576 net573 VPWR VGND sg13g2_buf_8
Xfanout562 net568 net562 VPWR VGND sg13g2_buf_8
Xfanout584 net591 net584 VPWR VGND sg13g2_buf_8
Xfanout595 _0639_ net595 VPWR VGND sg13g2_buf_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_34_619 VPWR VGND sg13g2_decap_4
XFILLER_26_181 VPWR VGND sg13g2_fill_2
XFILLER_10_571 VPWR VGND sg13g2_decap_4
XFILLER_6_542 VPWR VGND sg13g2_decap_4
XFILLER_6_586 VPWR VGND sg13g2_decap_8
XFILLER_6_564 VPWR VGND sg13g2_decap_4
XFILLER_29_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_240 VPWR VGND sg13g2_decap_8
X_4030_ _1744_ _1752_ _1753_ VPWR VGND sg13g2_nor2_1
XFILLER_46_991 VPWR VGND sg13g2_decap_8
X_4932_ net96 VGND VPWR _0483_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\]
+ _0140_ sg13g2_dfrbpq_1
XFILLER_24_129 VPWR VGND sg13g2_decap_8
X_4896__204 VPWR VGND net204 sg13g2_tiehi
X_4863_ net272 VGND VPWR _0414_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\]
+ _0071_ sg13g2_dfrbpq_1
X_4794_ net386 VGND VPWR _0345_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\]
+ _0045_ sg13g2_dfrbpq_1
X_3814_ net622 _1538_ _1543_ _1544_ VPWR VGND sg13g2_nor3_1
XFILLER_21_18 VPWR VGND sg13g2_fill_2
X_3745_ net596 VPWR _1475_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\]
+ net572 sg13g2_o21ai_1
X_4796__382 VPWR VGND net382 sg13g2_tiehi
X_4950__401 VPWR VGND net401 sg13g2_tiehi
X_3676_ net617 VPWR _1406_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\]
+ net586 sg13g2_o21ai_1
X_2627_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\] _0719_ _0591_
+ VPWR VGND sg13g2_mux2_1
X_2558_ _0673_ net600 _0672_ VPWR VGND sg13g2_nand2_2
X_4228_ _0875_ _0859_ _1935_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_424 VPWR VGND sg13g2_decap_8
XFILLER_29_925 VPWR VGND sg13g2_decap_8
X_4159_ _1866_ VPWR _1882_ VGND _1864_ _1881_ sg13g2_o21ai_1
XFILLER_28_446 VPWR VGND sg13g2_decap_8
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_23_140 VPWR VGND sg13g2_decap_8
XFILLER_24_674 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_fill_2
X_4938__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_7_339 VPWR VGND sg13g2_decap_8
XFILLER_3_523 VPWR VGND sg13g2_decap_8
XFILLER_11_84 VPWR VGND sg13g2_decap_8
XFILLER_47_711 VPWR VGND sg13g2_fill_1
XFILLER_35_928 VPWR VGND sg13g2_fill_2
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_28_991 VPWR VGND sg13g2_decap_8
X_5051__98 VPWR VGND net98 sg13g2_tiehi
X_3530_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\] net587 _1260_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_6_383 VPWR VGND sg13g2_decap_8
X_3461_ VGND VPWR _1191_ _1129_ net542 sg13g2_or2_1
X_3392_ _1122_ _1105_ _1107_ VPWR VGND sg13g2_xnor2_1
X_5062_ net240 VGND VPWR _0609_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\]
+ _0257_ sg13g2_dfrbpq_1
XFILLER_38_711 VPWR VGND sg13g2_fill_1
X_4013_ _1730_ _1643_ _1736_ VPWR VGND sg13g2_xor2_1
XFILLER_37_232 VPWR VGND sg13g2_fill_1
XFILLER_25_405 VPWR VGND sg13g2_fill_2
XFILLER_19_991 VPWR VGND sg13g2_decap_8
XFILLER_40_408 VPWR VGND sg13g2_decap_8
XFILLER_34_972 VPWR VGND sg13g2_decap_8
X_4915_ net166 VGND VPWR _0466_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\]
+ _0123_ sg13g2_dfrbpq_1
XFILLER_33_482 VPWR VGND sg13g2_decap_4
X_4846_ net305 VGND VPWR _0397_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[0\]
+ _0054_ sg13g2_dfrbpq_1
XFILLER_20_165 VPWR VGND sg13g2_decap_4
X_4777_ net48 VGND VPWR _0328_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\]
+ net634 sg13g2_dfrbpq_2
XFILLER_4_309 VPWR VGND sg13g2_fill_2
X_3728_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\] net579 _1458_ VPWR
+ VGND sg13g2_nor2_1
X_3659_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\] net584 _1389_ VPWR
+ VGND sg13g2_nor2_1
X_4718__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_0_548 VPWR VGND sg13g2_decap_8
XFILLER_28_210 VPWR VGND sg13g2_decap_8
XFILLER_17_928 VPWR VGND sg13g2_decap_8
XFILLER_28_276 VPWR VGND sg13g2_fill_2
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_32_909 VPWR VGND sg13g2_decap_8
XFILLER_25_983 VPWR VGND sg13g2_decap_8
XFILLER_8_604 VPWR VGND sg13g2_decap_8
XFILLER_8_637 VPWR VGND sg13g2_fill_2
XFILLER_12_688 VPWR VGND sg13g2_decap_4
XFILLER_11_198 VPWR VGND sg13g2_fill_1
XFILLER_4_887 VPWR VGND sg13g2_decap_8
XFILLER_35_714 VPWR VGND sg13g2_fill_2
XFILLER_47_585 VPWR VGND sg13g2_decap_8
XFILLER_16_950 VPWR VGND sg13g2_decap_8
X_2961_ VGND VPWR _0649_ net10 _0694_ _0671_ sg13g2_a21oi_2
XFILLER_31_920 VPWR VGND sg13g2_decap_8
XFILLER_34_268 VPWR VGND sg13g2_fill_1
X_4700_ net690 net744 _0253_ VPWR VGND sg13g2_nor2_1
X_2892_ _0725_ _0731_ _0783_ VPWR VGND sg13g2_nor2b_2
XFILLER_30_441 VPWR VGND sg13g2_fill_1
XFILLER_31_997 VPWR VGND sg13g2_decap_8
X_4631_ net688 net740 _0184_ VPWR VGND sg13g2_nor2_1
XFILLER_30_496 VPWR VGND sg13g2_decap_4
X_4562_ net681 net732 _0115_ VPWR VGND sg13g2_nor2_1
XFILLER_7_692 VPWR VGND sg13g2_decap_4
X_4493_ net651 net702 _0046_ VPWR VGND sg13g2_nor2_1
X_3513_ _1243_ _1158_ _1172_ VPWR VGND sg13g2_nand2_1
X_3444_ _1174_ _1004_ _1006_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_0 VPWR VGND sg13g2_decap_4
X_3375_ VPWR VGND _1103_ _1104_ _1073_ videogen.fancy_shader.n646\[7\] _1105_ net629
+ sg13g2_a221oi_1
X_5114_ net796 VGND VPWR serialize.n433\[1\] serialize.bit_cnt\[1\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_2
X_5045_ net181 VGND VPWR _0592_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\]
+ _0240_ sg13g2_dfrbpq_1
XFILLER_38_574 VPWR VGND sg13g2_decap_4
XFILLER_38_585 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_4
XFILLER_25_268 VPWR VGND sg13g2_fill_1
XFILLER_43_49 VPWR VGND sg13g2_fill_1
XFILLER_40_227 VPWR VGND sg13g2_decap_8
XFILLER_21_430 VPWR VGND sg13g2_fill_1
XFILLER_22_942 VPWR VGND sg13g2_decap_8
XFILLER_21_496 VPWR VGND sg13g2_fill_1
X_4829_ net330 VGND VPWR _0380_ tmds_red.n100 net649 sg13g2_dfrbpq_2
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_846 VPWR VGND sg13g2_decap_8
XFILLER_48_316 VPWR VGND sg13g2_decap_8
XFILLER_17_703 VPWR VGND sg13g2_fill_1
XFILLER_44_511 VPWR VGND sg13g2_fill_1
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_566 VPWR VGND sg13g2_decap_8
XFILLER_16_235 VPWR VGND sg13g2_fill_1
XFILLER_17_769 VPWR VGND sg13g2_fill_1
XFILLER_44_599 VPWR VGND sg13g2_decap_4
XFILLER_44_577 VPWR VGND sg13g2_fill_1
XFILLER_16_279 VPWR VGND sg13g2_fill_2
XFILLER_8_401 VPWR VGND sg13g2_decap_8
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_12_441 VPWR VGND sg13g2_fill_1
XFILLER_12_452 VPWR VGND sg13g2_decap_8
XFILLER_13_986 VPWR VGND sg13g2_decap_8
XFILLER_33_82 VPWR VGND sg13g2_fill_1
XFILLER_8_489 VPWR VGND sg13g2_decap_8
XFILLER_8_478 VPWR VGND sg13g2_fill_2
XFILLER_3_161 VPWR VGND sg13g2_fill_1
XFILLER_3_194 VPWR VGND sg13g2_fill_1
X_3160_ _0929_ VPWR _0930_ VGND videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ _0928_ sg13g2_o21ai_1
XFILLER_12_4 VPWR VGND sg13g2_fill_1
X_3091_ _0878_ _0880_ _0881_ VPWR VGND sg13g2_nor2_1
Xhold1 clockdiv.q2 VPWR VGND net406 sg13g2_dlygate4sd3_1
XFILLER_35_533 VPWR VGND sg13g2_decap_8
XFILLER_35_577 VPWR VGND sg13g2_fill_2
XFILLER_35_599 VPWR VGND sg13g2_decap_8
X_3993_ _1548_ _1352_ _1718_ _1719_ VPWR VGND sg13g2_a21o_1
X_2944_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0792_ _0802_ VPWR
+ VGND sg13g2_and2_1
X_2875_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\] net772 _0779_ _0394_
+ VPWR VGND sg13g2_mux2_1
X_4614_ net691 net743 _0167_ VPWR VGND sg13g2_nor2_1
X_4545_ net661 net712 _0098_ VPWR VGND sg13g2_nor2_1
X_4476_ net653 net704 _0029_ VPWR VGND sg13g2_nor2_1
X_3427_ _1153_ _1155_ _1036_ _1157_ VPWR VGND sg13g2_nand3_1
X_3358_ _1088_ _1087_ VPWR VGND sg13g2_inv_2
XFILLER_39_861 VPWR VGND sg13g2_decap_8
X_3289_ _1019_ _1010_ _1018_ VPWR VGND sg13g2_nand2_1
X_5028_ net318 VGND VPWR _0575_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\]
+ _0223_ sg13g2_dfrbpq_1
XFILLER_26_522 VPWR VGND sg13g2_decap_8
XFILLER_13_249 VPWR VGND sg13g2_decap_4
XFILLER_10_912 VPWR VGND sg13g2_decap_8
XFILLER_22_761 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_10_989 VPWR VGND sg13g2_decap_8
X_4747__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_1_676 VPWR VGND sg13g2_decap_8
XFILLER_1_687 VPWR VGND sg13g2_fill_2
XFILLER_23_1018 VPWR VGND sg13g2_decap_8
XFILLER_28_93 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_decap_8
XFILLER_44_396 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_fill_1
XFILLER_8_220 VPWR VGND sg13g2_decap_8
XFILLER_9_721 VPWR VGND sg13g2_decap_8
XFILLER_8_231 VPWR VGND sg13g2_fill_2
X_2660_ _0679_ _0712_ _0731_ VPWR VGND sg13g2_nor2_2
XFILLER_5_960 VPWR VGND sg13g2_decap_8
X_2591_ net588 _0701_ _0702_ VPWR VGND sg13g2_nor2_2
XFILLER_4_470 VPWR VGND sg13g2_decap_4
X_4330_ _2026_ net602 _2023_ VPWR VGND sg13g2_nand2_1
X_4261_ _1965_ _1966_ _1967_ VPWR VGND sg13g2_and2_1
X_3212_ net751 _0963_ _0349_ VPWR VGND sg13g2_nor2_1
X_4192_ _1900_ VPWR _1911_ VGND _1902_ _1904_ sg13g2_o21ai_1
X_3143_ _0918_ _0665_ _0670_ VPWR VGND sg13g2_nand2_2
X_3074_ _0864_ tmds_red.n102 _0862_ VPWR VGND sg13g2_nand2_1
XFILLER_39_1014 VPWR VGND sg13g2_decap_8
XFILLER_36_886 VPWR VGND sg13g2_fill_2
XFILLER_23_536 VPWR VGND sg13g2_fill_1
X_4979__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_11_709 VPWR VGND sg13g2_decap_4
XFILLER_23_569 VPWR VGND sg13g2_decap_8
X_3976_ _1625_ _1701_ _1702_ VPWR VGND sg13g2_nor2_1
X_2927_ _0790_ _0715_ _0763_ VPWR VGND sg13g2_nand2_2
X_2858_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\] net756 _0776_ _0408_
+ VPWR VGND sg13g2_mux2_1
X_2789_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\] net767 _0758_ _0459_
+ VPWR VGND sg13g2_mux2_1
X_4528_ net657 net708 _0081_ VPWR VGND sg13g2_nor2_1
XFILLER_2_407 VPWR VGND sg13g2_decap_8
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_1
X_4459_ net656 net702 _0012_ VPWR VGND sg13g2_nor2_1
Xfanout722 net723 net722 VPWR VGND sg13g2_buf_8
Xfanout733 net734 net733 VPWR VGND sg13g2_buf_8
Xfanout711 net746 net711 VPWR VGND sg13g2_buf_8
Xfanout744 net745 net744 VPWR VGND sg13g2_buf_8
Xfanout755 net761 net755 VPWR VGND sg13g2_buf_8
Xfanout766 ui_in[6] net766 VPWR VGND sg13g2_buf_8
Xfanout799 net802 net799 VPWR VGND sg13g2_buf_8
Xfanout788 net791 net788 VPWR VGND sg13g2_buf_8
Xfanout777 net781 net777 VPWR VGND sg13g2_buf_8
XFILLER_39_680 VPWR VGND sg13g2_fill_1
XFILLER_14_525 VPWR VGND sg13g2_decap_8
X_4993__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_14_73 VPWR VGND sg13g2_fill_1
XFILLER_5_267 VPWR VGND sg13g2_fill_1
XFILLER_2_930 VPWR VGND sg13g2_decap_8
XFILLER_49_433 VPWR VGND sg13g2_decap_8
XFILLER_1_495 VPWR VGND sg13g2_fill_2
XFILLER_49_455 VPWR VGND sg13g2_decap_8
XFILLER_33_845 VPWR VGND sg13g2_decap_8
X_3830_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\] net566 _1559_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_366 VPWR VGND sg13g2_decap_8
XFILLER_33_878 VPWR VGND sg13g2_fill_2
X_3761_ net599 VPWR _1491_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\]
+ net552 sg13g2_o21ai_1
XFILLER_20_528 VPWR VGND sg13g2_decap_4
X_2712_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\] _0742_ _0529_
+ VPWR VGND sg13g2_mux2_1
X_3692_ net592 _1416_ _1421_ _1422_ VPWR VGND sg13g2_nor3_1
X_2643_ _0714_ _0725_ _0726_ VPWR VGND sg13g2_nor2_2
X_2574_ _0689_ _0680_ VPWR VGND _0687_ sg13g2_nand2b_2
X_4313_ VGND VPWR _2010_ _2012_ _0616_ net749 sg13g2_a21oi_1
X_4244_ _0889_ _1950_ _1951_ VPWR VGND sg13g2_nor2_1
X_4175_ _1895_ VPWR _1898_ VGND _1896_ _1897_ sg13g2_o21ai_1
X_4866__267 VPWR VGND net267 sg13g2_tiehi
X_3126_ _0800_ _0898_ _0905_ _0309_ VPWR VGND sg13g2_nor3_1
X_3057_ _0847_ tmds_green.n126 _0848_ VPWR VGND sg13g2_xor2_1
XFILLER_11_517 VPWR VGND sg13g2_decap_8
X_3959_ _1671_ _1682_ _1629_ _1685_ VPWR VGND sg13g2_nand3_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_4873__249 VPWR VGND net249 sg13g2_tiehi
XFILLER_3_716 VPWR VGND sg13g2_decap_8
XFILLER_2_204 VPWR VGND sg13g2_decap_8
Xfanout563 net564 net563 VPWR VGND sg13g2_buf_8
Xfanout552 net558 net552 VPWR VGND sg13g2_buf_8
Xfanout574 net576 net574 VPWR VGND sg13g2_buf_8
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_46_425 VPWR VGND sg13g2_decap_8
X_4845__307 VPWR VGND net307 sg13g2_tiehi
XFILLER_18_105 VPWR VGND sg13g2_fill_1
Xfanout596 net599 net596 VPWR VGND sg13g2_buf_8
Xfanout585 net591 net585 VPWR VGND sg13g2_buf_8
XFILLER_15_812 VPWR VGND sg13g2_decap_8
XFILLER_27_661 VPWR VGND sg13g2_decap_4
XFILLER_42_631 VPWR VGND sg13g2_fill_1
XFILLER_14_311 VPWR VGND sg13g2_decap_8
XFILLER_15_823 VPWR VGND sg13g2_fill_1
XFILLER_26_171 VPWR VGND sg13g2_decap_4
XFILLER_41_141 VPWR VGND sg13g2_decap_8
XFILLER_14_355 VPWR VGND sg13g2_decap_4
XFILLER_15_856 VPWR VGND sg13g2_fill_1
XFILLER_30_859 VPWR VGND sg13g2_decap_4
XFILLER_6_554 VPWR VGND sg13g2_decap_4
XFILLER_6_532 VPWR VGND sg13g2_fill_1
XFILLER_29_1002 VPWR VGND sg13g2_decap_8
XFILLER_1_281 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_38_926 VPWR VGND sg13g2_fill_1
XFILLER_49_296 VPWR VGND sg13g2_decap_8
XFILLER_37_447 VPWR VGND sg13g2_fill_1
XFILLER_2_87 VPWR VGND sg13g2_decap_4
XFILLER_46_970 VPWR VGND sg13g2_decap_8
XFILLER_25_609 VPWR VGND sg13g2_fill_2
XFILLER_45_491 VPWR VGND sg13g2_decap_4
X_4931_ net100 VGND VPWR _0482_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\]
+ _0139_ sg13g2_dfrbpq_1
X_4862_ net274 VGND VPWR _0413_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\]
+ _0070_ sg13g2_dfrbpq_1
XFILLER_21_804 VPWR VGND sg13g2_fill_1
X_3813_ _1539_ _1540_ _1541_ _1542_ _1543_ VPWR VGND sg13g2_nor4_1
X_4793_ net388 VGND VPWR _0344_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\]
+ _0044_ sg13g2_dfrbpq_1
X_3744_ net613 VPWR _1474_ VGND _1467_ _1473_ sg13g2_o21ai_1
X_3675_ _1401_ _1402_ _1403_ _1404_ _1405_ VPWR VGND sg13g2_nor4_1
X_2626_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\] _0719_ _0592_
+ VPWR VGND sg13g2_mux2_1
X_2557_ _0665_ _0671_ _0672_ VPWR VGND sg13g2_nor2_2
X_4227_ tmds_red.dc_balancing_reg\[1\] _0859_ _1934_ VPWR VGND sg13g2_nor2_1
XFILLER_29_904 VPWR VGND sg13g2_decap_8
X_4983__266 VPWR VGND net266 sg13g2_tiehi
X_4158_ VGND VPWR _1866_ _1869_ _1881_ _1860_ sg13g2_a21oi_1
XFILLER_44_918 VPWR VGND sg13g2_decap_8
X_4089_ _1804_ _1084_ _1812_ VPWR VGND sg13g2_xor2_1
X_3109_ net569 _0895_ _0278_ VPWR VGND sg13g2_nor2_1
XFILLER_24_642 VPWR VGND sg13g2_decap_4
XFILLER_11_303 VPWR VGND sg13g2_decap_8
XFILLER_11_314 VPWR VGND sg13g2_fill_2
XFILLER_23_163 VPWR VGND sg13g2_fill_1
XFILLER_3_502 VPWR VGND sg13g2_fill_1
XFILLER_46_244 VPWR VGND sg13g2_decap_8
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_fill_2
XFILLER_43_984 VPWR VGND sg13g2_decap_8
XFILLER_14_174 VPWR VGND sg13g2_decap_4
XFILLER_7_852 VPWR VGND sg13g2_decap_8
XFILLER_7_830 VPWR VGND sg13g2_fill_1
XFILLER_11_881 VPWR VGND sg13g2_decap_4
X_3460_ net542 _1129_ _1088_ _1190_ VPWR VGND sg13g2_nand3_1
XFILLER_6_373 VPWR VGND sg13g2_decap_4
X_3391_ VPWR _1121_ _1120_ VGND sg13g2_inv_1
X_5061_ net260 VGND VPWR _0608_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\]
+ _0256_ sg13g2_dfrbpq_1
XFILLER_42_1021 VPWR VGND sg13g2_decap_8
X_4012_ _1733_ _1734_ _1735_ VPWR VGND sg13g2_and2_1
XFILLER_19_970 VPWR VGND sg13g2_decap_8
XFILLER_18_480 VPWR VGND sg13g2_fill_2
X_4914_ net168 VGND VPWR _0465_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\]
+ _0122_ sg13g2_dfrbpq_1
X_4845_ net307 VGND VPWR _0396_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\]
+ _0053_ sg13g2_dfrbpq_1
XFILLER_20_122 VPWR VGND sg13g2_decap_8
XFILLER_21_645 VPWR VGND sg13g2_decap_8
X_4776_ net50 VGND VPWR _0327_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\]
+ net632 sg13g2_dfrbpq_2
X_3727_ net598 VPWR _1457_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\]
+ net555 sg13g2_o21ai_1
X_3658_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\] net574 _1388_ VPWR
+ VGND sg13g2_nor2_1
X_2609_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\] _0711_ _0601_
+ VPWR VGND sg13g2_mux2_1
X_3589_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\] net574 _1319_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_48_509 VPWR VGND sg13g2_fill_1
X_4909__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_44_748 VPWR VGND sg13g2_fill_1
XFILLER_44_759 VPWR VGND sg13g2_decap_4
XFILLER_25_962 VPWR VGND sg13g2_decap_8
XFILLER_12_601 VPWR VGND sg13g2_decap_8
XFILLER_19_1012 VPWR VGND sg13g2_decap_8
XFILLER_19_1023 VPWR VGND sg13g2_fill_2
XFILLER_40_998 VPWR VGND sg13g2_decap_8
XFILLER_8_627 VPWR VGND sg13g2_fill_2
XFILLER_4_800 VPWR VGND sg13g2_fill_1
XFILLER_3_354 VPWR VGND sg13g2_fill_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_47_564 VPWR VGND sg13g2_decap_8
XFILLER_34_247 VPWR VGND sg13g2_decap_8
XFILLER_43_781 VPWR VGND sg13g2_fill_2
X_2960_ VGND VPWR _0649_ net9 _0691_ _0671_ sg13g2_a21oi_2
X_2891_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\] _0782_ _0338_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_20 VPWR VGND sg13g2_decap_4
X_4630_ net692 net740 _0183_ VPWR VGND sg13g2_nor2_1
XFILLER_31_976 VPWR VGND sg13g2_decap_8
X_4561_ net681 net732 _0114_ VPWR VGND sg13g2_nor2_1
X_4492_ net652 net703 _0045_ VPWR VGND sg13g2_nor2_1
X_3512_ VPWR VGND _1186_ net547 _1179_ net545 _1242_ _1170_ sg13g2_a221oi_1
XFILLER_6_181 VPWR VGND sg13g2_fill_2
X_3443_ _1173_ _1171_ _1172_ VPWR VGND sg13g2_nand2_1
X_5113_ net796 VGND VPWR serialize.n433\[0\] serialize.bit_cnt\[0\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_2
X_3374_ _1074_ _1101_ _1104_ VPWR VGND sg13g2_nor2_1
XFILLER_33_0 VPWR VGND sg13g2_decap_8
X_5044_ net189 VGND VPWR _0591_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\]
+ _0239_ sg13g2_dfrbpq_1
XFILLER_22_921 VPWR VGND sg13g2_decap_8
XFILLER_21_442 VPWR VGND sg13g2_decap_8
X_4828_ net331 VGND VPWR _0379_ tmds_red.n102 net644 sg13g2_dfrbpq_2
X_4774__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_22_998 VPWR VGND sg13g2_decap_8
X_4759_ net80 VGND VPWR _0310_ videogen.fancy_shader.video_x\[7\] net638 sg13g2_dfrbpq_1
XFILLER_49_1016 VPWR VGND sg13g2_decap_8
XFILLER_49_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_825 VPWR VGND sg13g2_decap_8
XFILLER_0_379 VPWR VGND sg13g2_decap_8
XFILLER_1_1007 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_decap_4
XFILLER_16_203 VPWR VGND sg13g2_decap_8
XFILLER_29_586 VPWR VGND sg13g2_decap_8
XFILLER_16_258 VPWR VGND sg13g2_decap_8
XFILLER_17_95 VPWR VGND sg13g2_fill_2
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_25_781 VPWR VGND sg13g2_decap_4
XFILLER_31_228 VPWR VGND sg13g2_decap_8
XFILLER_13_965 VPWR VGND sg13g2_decap_8
XFILLER_12_475 VPWR VGND sg13g2_fill_2
XFILLER_33_72 VPWR VGND sg13g2_decap_4
XFILLER_4_630 VPWR VGND sg13g2_decap_4
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_0_891 VPWR VGND sg13g2_decap_8
X_3090_ _0880_ _0879_ VPWR VGND sg13g2_inv_2
Xhold2 _0623_ VPWR VGND net407 sg13g2_dlygate4sd3_1
XFILLER_48_895 VPWR VGND sg13g2_decap_8
XFILLER_47_372 VPWR VGND sg13g2_decap_8
XFILLER_35_512 VPWR VGND sg13g2_fill_2
XFILLER_22_206 VPWR VGND sg13g2_fill_1
X_3992_ _1451_ VPWR _1718_ VGND _1352_ _1548_ sg13g2_o21ai_1
X_2943_ net629 _0666_ _0801_ VPWR VGND sg13g2_nor2b_1
X_2874_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\] net762 _0779_ _0395_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_773 VPWR VGND sg13g2_decap_8
X_4613_ net690 net744 _0166_ VPWR VGND sg13g2_nor2_1
X_4544_ net679 net730 _0097_ VPWR VGND sg13g2_nor2_1
X_4475_ net668 net720 _0028_ VPWR VGND sg13g2_nor2_1
X_3426_ VGND VPWR _1153_ _1155_ _1156_ _1036_ sg13g2_a21oi_1
X_3357_ _1085_ _1086_ _1087_ VPWR VGND sg13g2_and2_1
X_5027_ net349 VGND VPWR _0574_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\]
+ _0222_ sg13g2_dfrbpq_1
X_3288_ _1016_ _1014_ _1018_ VPWR VGND sg13g2_xor2_1
X_5045__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_41_537 VPWR VGND sg13g2_fill_2
XFILLER_21_250 VPWR VGND sg13g2_fill_1
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_10_968 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_fill_2
XFILLER_5_416 VPWR VGND sg13g2_decap_8
XFILLER_49_637 VPWR VGND sg13g2_decap_8
XFILLER_0_198 VPWR VGND sg13g2_fill_2
XFILLER_28_50 VPWR VGND sg13g2_decap_4
XFILLER_45_887 VPWR VGND sg13g2_decap_8
XFILLER_32_548 VPWR VGND sg13g2_fill_1
XFILLER_13_762 VPWR VGND sg13g2_decap_8
XFILLER_13_784 VPWR VGND sg13g2_fill_1
XFILLER_13_795 VPWR VGND sg13g2_decap_4
XFILLER_9_755 VPWR VGND sg13g2_fill_2
XFILLER_9_788 VPWR VGND sg13g2_decap_8
XFILLER_9_799 VPWR VGND sg13g2_fill_1
X_2590_ _0701_ net600 _0695_ VPWR VGND sg13g2_nand2_2
XFILLER_5_87 VPWR VGND sg13g2_fill_1
XFILLER_5_65 VPWR VGND sg13g2_fill_1
X_4260_ VGND VPWR _1933_ _1941_ _1966_ _1943_ sg13g2_a21oi_1
X_3211_ _0963_ videogen.fancy_shader.n646\[3\] _0961_ VPWR VGND sg13g2_xnor2_1
X_4191_ _1910_ VPWR _0382_ VGND net750 _1909_ sg13g2_o21ai_1
X_3142_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0916_ _0917_ VPWR VGND
+ sg13g2_nor2_1
XFILLER_39_158 VPWR VGND sg13g2_decap_8
X_3073_ tmds_red.n102 _0862_ _0863_ VPWR VGND sg13g2_nor2_1
XFILLER_23_548 VPWR VGND sg13g2_decap_8
X_3975_ _1700_ _1699_ _1234_ _1701_ VPWR VGND sg13g2_a21o_1
X_2926_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\] net783 _0789_ _0279_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_581 VPWR VGND sg13g2_fill_2
X_2857_ _0718_ _0772_ _0776_ VPWR VGND sg13g2_nor2_2
X_2788_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\] net757 _0758_ _0460_
+ VPWR VGND sg13g2_mux2_1
X_4527_ net658 net709 _0080_ VPWR VGND sg13g2_nor2_1
XFILLER_46_1019 VPWR VGND sg13g2_decap_8
X_4458_ net651 net707 _0011_ VPWR VGND sg13g2_nor2_1
XFILLER_49_49 VPWR VGND sg13g2_decap_8
Xfanout701 serialize.n410 net701 VPWR VGND sg13g2_buf_2
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_2
X_3409_ _1121_ VPWR _1139_ VGND _1115_ _1137_ sg13g2_o21ai_1
Xfanout712 net714 net712 VPWR VGND sg13g2_buf_8
X_4389_ _2076_ _2079_ _2080_ VPWR VGND sg13g2_nor2_2
Xfanout767 net768 net767 VPWR VGND sg13g2_buf_8
Xfanout734 net746 net734 VPWR VGND sg13g2_buf_8
Xfanout756 net760 net756 VPWR VGND sg13g2_buf_8
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
Xfanout778 net781 net778 VPWR VGND sg13g2_buf_8
Xfanout789 net791 net789 VPWR VGND sg13g2_buf_8
XFILLER_26_353 VPWR VGND sg13g2_decap_8
XFILLER_26_364 VPWR VGND sg13g2_fill_1
XFILLER_27_898 VPWR VGND sg13g2_decap_8
XFILLER_6_714 VPWR VGND sg13g2_decap_8
XFILLER_49_401 VPWR VGND sg13g2_decap_8
XFILLER_7_1024 VPWR VGND sg13g2_decap_4
XFILLER_2_986 VPWR VGND sg13g2_decap_8
X_4965__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_37_618 VPWR VGND sg13g2_fill_2
XFILLER_18_832 VPWR VGND sg13g2_decap_8
XFILLER_44_150 VPWR VGND sg13g2_decap_4
XFILLER_18_876 VPWR VGND sg13g2_decap_8
XFILLER_33_813 VPWR VGND sg13g2_decap_4
XFILLER_17_397 VPWR VGND sg13g2_fill_1
XFILLER_44_194 VPWR VGND sg13g2_fill_2
X_3760_ _1486_ _1487_ _1488_ _1489_ _1490_ VPWR VGND sg13g2_nor4_1
XFILLER_20_507 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_fill_1
X_4972__308 VPWR VGND net308 sg13g2_tiehi
X_2711_ _0742_ _0706_ _0717_ VPWR VGND sg13g2_nand2_2
XFILLER_9_574 VPWR VGND sg13g2_decap_4
X_3691_ _1417_ _1418_ _1419_ _1420_ _1421_ VPWR VGND sg13g2_nor4_1
X_2642_ _0692_ _0697_ net619 _0725_ VPWR VGND sg13g2_nand3_1
X_2573_ _0679_ _0687_ _0688_ VPWR VGND sg13g2_nor2_2
X_4312_ _1999_ _2011_ _2012_ VPWR VGND sg13g2_nor2_1
X_4243_ VGND VPWR _0855_ _1929_ _1950_ _1939_ sg13g2_a21oi_1
XFILLER_19_19 VPWR VGND sg13g2_fill_1
X_4174_ _1897_ net547 _1235_ VPWR VGND sg13g2_nand2_1
X_3125_ videogen.fancy_shader.video_x\[6\] _0799_ _0905_ VPWR VGND sg13g2_nor2_1
XFILLER_27_106 VPWR VGND sg13g2_fill_1
X_3056_ _0846_ VPWR _0847_ VGND _0839_ _0843_ sg13g2_o21ai_1
XFILLER_24_835 VPWR VGND sg13g2_decap_8
XFILLER_23_334 VPWR VGND sg13g2_decap_8
XFILLER_23_378 VPWR VGND sg13g2_decap_8
XFILLER_13_1007 VPWR VGND sg13g2_decap_8
X_3958_ _1683_ _1671_ _1629_ _1684_ VPWR VGND sg13g2_a21o_1
X_3889_ VGND VPWR net1 _1250_ _1618_ _1617_ sg13g2_a21oi_1
X_2909_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\] _0786_ _0293_
+ VPWR VGND sg13g2_mux2_1
Xfanout542 _1111_ net542 VPWR VGND sg13g2_buf_8
Xfanout553 net557 net553 VPWR VGND sg13g2_buf_8
Xfanout564 net567 net564 VPWR VGND sg13g2_buf_8
Xfanout575 net576 net575 VPWR VGND sg13g2_buf_8
XFILLER_47_927 VPWR VGND sg13g2_decap_8
Xfanout586 net590 net586 VPWR VGND sg13g2_buf_8
Xfanout597 net599 net597 VPWR VGND sg13g2_buf_8
XFILLER_42_654 VPWR VGND sg13g2_decap_4
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_25_51 VPWR VGND sg13g2_decap_4
XFILLER_26_194 VPWR VGND sg13g2_decap_4
XFILLER_25_84 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_fill_1
XFILLER_30_827 VPWR VGND sg13g2_fill_2
X_4919__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_41_83 VPWR VGND sg13g2_decap_4
XFILLER_37_7 VPWR VGND sg13g2_fill_1
XFILLER_2_794 VPWR VGND sg13g2_decap_8
XFILLER_18_640 VPWR VGND sg13g2_fill_2
XFILLER_18_651 VPWR VGND sg13g2_fill_1
X_4930_ net104 VGND VPWR _0481_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\]
+ _0138_ sg13g2_dfrbpq_1
X_4861_ net276 VGND VPWR _0412_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\]
+ _0069_ sg13g2_dfrbpq_1
X_3812_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\] net566 _1542_ VPWR
+ VGND sg13g2_nor2_1
X_4792_ net390 VGND VPWR _0343_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\]
+ _0043_ sg13g2_dfrbpq_1
XFILLER_21_849 VPWR VGND sg13g2_fill_2
X_3743_ net620 VPWR _1473_ VGND _1468_ _1472_ sg13g2_o21ai_1
X_3674_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\] net587 _1404_ VPWR
+ VGND sg13g2_nor2_1
X_2625_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\] _0719_ _0593_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_709 VPWR VGND sg13g2_decap_8
X_2556_ _0668_ _0669_ _0667_ _0671_ VPWR VGND sg13g2_nand3_1
X_4226_ VPWR _1933_ _1932_ VGND sg13g2_inv_1
X_4157_ _1876_ _1879_ _1880_ VPWR VGND sg13g2_nor2_1
X_3108_ _0895_ _0854_ _0894_ VPWR VGND sg13g2_xnor2_1
X_4088_ _1811_ _1124_ _1809_ VPWR VGND sg13g2_xnor2_1
X_3039_ _0807_ _0810_ _0000_ VPWR VGND sg13g2_nor2_1
XFILLER_11_337 VPWR VGND sg13g2_decap_8
XFILLER_11_348 VPWR VGND sg13g2_fill_2
XFILLER_20_860 VPWR VGND sg13g2_fill_1
XFILLER_11_64 VPWR VGND sg13g2_fill_2
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_415 VPWR VGND sg13g2_decap_4
XFILLER_46_267 VPWR VGND sg13g2_decap_8
XFILLER_46_278 VPWR VGND sg13g2_fill_1
XFILLER_34_429 VPWR VGND sg13g2_fill_1
XFILLER_43_963 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_6_330 VPWR VGND sg13g2_decap_4
X_3390_ _1120_ _1117_ _1119_ VPWR VGND sg13g2_xnor2_1
X_5060_ net275 VGND VPWR _0607_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\]
+ _0255_ sg13g2_dfrbpq_1
XFILLER_42_1000 VPWR VGND sg13g2_decap_8
X_4011_ _1734_ _1731_ _1732_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_919 VPWR VGND sg13g2_decap_8
X_4913_ net170 VGND VPWR _0464_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[3\]
+ _0121_ sg13g2_dfrbpq_1
XFILLER_33_451 VPWR VGND sg13g2_decap_4
X_4844_ net309 VGND VPWR _0395_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\]
+ _0052_ sg13g2_dfrbpq_1
X_4775_ net52 VGND VPWR _0326_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\]
+ net634 sg13g2_dfrbpq_1
XFILLER_21_657 VPWR VGND sg13g2_fill_2
X_3726_ _1452_ _1453_ _1454_ _1455_ _1456_ VPWR VGND sg13g2_nor4_1
X_3657_ net615 VPWR _1387_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\]
+ net552 sg13g2_o21ai_1
X_2608_ _0711_ _0688_ _0710_ VPWR VGND sg13g2_nand2_2
X_3588_ net620 VPWR _1318_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\]
+ net585 sg13g2_o21ai_1
X_2539_ VPWR _0656_ net414 VGND sg13g2_inv_1
XFILLER_29_724 VPWR VGND sg13g2_decap_4
X_4209_ net751 _1923_ _0387_ VPWR VGND sg13g2_nor2_1
XFILLER_25_941 VPWR VGND sg13g2_decap_8
XFILLER_40_900 VPWR VGND sg13g2_decap_4
XFILLER_12_624 VPWR VGND sg13g2_decap_8
XFILLER_40_977 VPWR VGND sg13g2_decap_8
XFILLER_11_134 VPWR VGND sg13g2_fill_1
XFILLER_11_145 VPWR VGND sg13g2_fill_2
XFILLER_8_639 VPWR VGND sg13g2_fill_1
XFILLER_22_52 VPWR VGND sg13g2_decap_8
XFILLER_7_149 VPWR VGND sg13g2_decap_8
XFILLER_22_85 VPWR VGND sg13g2_decap_8
XFILLER_3_311 VPWR VGND sg13g2_fill_2
XFILLER_22_96 VPWR VGND sg13g2_fill_2
XFILLER_3_366 VPWR VGND sg13g2_decap_8
XFILLER_26_1017 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_28_790 VPWR VGND sg13g2_fill_1
XFILLER_16_985 VPWR VGND sg13g2_decap_8
XFILLER_30_410 VPWR VGND sg13g2_decap_8
X_2890_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\] _0782_ _0339_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_955 VPWR VGND sg13g2_decap_8
XFILLER_30_454 VPWR VGND sg13g2_decap_4
XFILLER_8_43 VPWR VGND sg13g2_fill_1
X_4560_ net681 net732 _0113_ VPWR VGND sg13g2_nor2_1
X_4491_ net653 net704 _0044_ VPWR VGND sg13g2_nor2_1
X_3511_ _1188_ _1189_ _1179_ _1241_ VPWR VGND _1240_ sg13g2_nand4_1
X_3442_ _1022_ VPWR _1172_ VGND _1165_ _1169_ sg13g2_o21ai_1
X_3373_ _1075_ _1102_ _1103_ VPWR VGND sg13g2_nor2_1
X_5112_ net797 VGND VPWR serialize.n429\[9\] serialize.n417\[7\] clknet_3_0__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
X_5043_ net197 VGND VPWR _0590_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\]
+ _0238_ sg13g2_dfrbpq_1
XFILLER_27_19 VPWR VGND sg13g2_decap_8
XFILLER_26_738 VPWR VGND sg13g2_fill_1
XFILLER_26_749 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_25_259 VPWR VGND sg13g2_fill_2
XFILLER_21_410 VPWR VGND sg13g2_decap_8
XFILLER_22_977 VPWR VGND sg13g2_decap_8
X_4827_ net332 VGND VPWR _0378_ tmds_green.n132 net647 sg13g2_dfrbpq_1
XFILLER_21_476 VPWR VGND sg13g2_fill_2
X_4758_ net81 VGND VPWR _0309_ videogen.fancy_shader.video_x\[6\] net638 sg13g2_dfrbpq_2
X_4689_ net686 net737 _0242_ VPWR VGND sg13g2_nor2_1
X_3709_ _1435_ _1436_ _1437_ _1438_ _1439_ VPWR VGND sg13g2_nor4_1
XFILLER_1_804 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_48_307 VPWR VGND sg13g2_decap_4
XFILLER_44_502 VPWR VGND sg13g2_decap_8
XFILLER_17_716 VPWR VGND sg13g2_decap_8
XFILLER_44_546 VPWR VGND sg13g2_fill_2
XFILLER_44_535 VPWR VGND sg13g2_decap_8
X_4996__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_32_708 VPWR VGND sg13g2_decap_8
XFILLER_13_944 VPWR VGND sg13g2_decap_8
XFILLER_12_432 VPWR VGND sg13g2_decap_8
XFILLER_8_436 VPWR VGND sg13g2_fill_2
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_8_447 VPWR VGND sg13g2_fill_1
XFILLER_4_675 VPWR VGND sg13g2_decap_8
Xhold3 serialize.n420\[1\] VPWR VGND net408 sg13g2_dlygate4sd3_1
XFILLER_0_870 VPWR VGND sg13g2_decap_8
XFILLER_48_874 VPWR VGND sg13g2_decap_8
X_3991_ _1352_ _1548_ _1717_ VPWR VGND sg13g2_nor2_1
XFILLER_35_579 VPWR VGND sg13g2_fill_1
X_2942_ videogen.fancy_shader.video_x\[6\] _0799_ _0800_ VPWR VGND sg13g2_and2_1
X_2873_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\] net752 _0779_ _0396_
+ VPWR VGND sg13g2_mux2_1
X_4612_ net692 net744 _0165_ VPWR VGND sg13g2_nor2_1
X_4801__372 VPWR VGND net372 sg13g2_tiehi
XFILLER_30_284 VPWR VGND sg13g2_fill_2
X_4543_ net680 net731 _0096_ VPWR VGND sg13g2_nor2_1
X_4474_ net659 net710 _0027_ VPWR VGND sg13g2_nor2_1
X_3425_ _1140_ _1136_ _1154_ _1155_ VPWR VGND sg13g2_a21o_2
X_3356_ _1086_ _1076_ _1084_ VPWR VGND sg13g2_nand2b_1
X_3287_ _1017_ _1014_ _1016_ VPWR VGND sg13g2_nand2b_1
X_5026_ net357 VGND VPWR _0573_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\]
+ _0221_ sg13g2_dfrbpq_1
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_22_796 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_10_947 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_48_115 VPWR VGND sg13g2_fill_2
XFILLER_0_177 VPWR VGND sg13g2_decap_8
XFILLER_29_351 VPWR VGND sg13g2_decap_4
XFILLER_44_310 VPWR VGND sg13g2_fill_1
XFILLER_17_535 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_fill_1
XFILLER_44_365 VPWR VGND sg13g2_decap_8
XFILLER_44_376 VPWR VGND sg13g2_fill_1
XFILLER_5_995 VPWR VGND sg13g2_decap_8
X_3210_ _0961_ _0962_ _0348_ VPWR VGND sg13g2_nor2_1
X_4190_ _1910_ _1616_ _1905_ VPWR VGND sg13g2_nand2_1
X_3141_ _0913_ _0915_ _0916_ VPWR VGND sg13g2_nor2b_1
X_3072_ _0862_ _0859_ _0861_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_505 VPWR VGND sg13g2_fill_2
XFILLER_35_365 VPWR VGND sg13g2_decap_8
XFILLER_35_376 VPWR VGND sg13g2_fill_1
X_3974_ VGND VPWR _1700_ _1698_ _1686_ sg13g2_or2_1
X_2925_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[1\] net772 _0789_ _0280_
+ VPWR VGND sg13g2_mux2_1
X_2856_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\] _0775_ _0409_
+ VPWR VGND sg13g2_mux2_1
XFILLER_40_19 VPWR VGND sg13g2_decap_8
X_2787_ _0725_ _0751_ _0758_ VPWR VGND sg13g2_nor2b_2
X_4526_ net657 net708 _0079_ VPWR VGND sg13g2_nor2_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
X_4457_ net657 net708 _0010_ VPWR VGND sg13g2_nor2_1
X_3408_ _1120_ _1126_ _1138_ VPWR VGND _1137_ sg13g2_nand3b_1
Xfanout702 net703 net702 VPWR VGND sg13g2_buf_8
Xfanout724 net746 net724 VPWR VGND sg13g2_buf_8
Xfanout713 net714 net713 VPWR VGND sg13g2_buf_1
X_4388_ VGND VPWR _1995_ _2077_ _2079_ _2078_ sg13g2_a21oi_1
Xfanout757 net760 net757 VPWR VGND sg13g2_buf_8
Xfanout746 clockdiv.q1 net746 VPWR VGND sg13g2_buf_8
Xfanout735 net739 net735 VPWR VGND sg13g2_buf_8
X_3339_ VPWR _1069_ _1068_ VGND sg13g2_inv_1
Xfanout768 net771 net768 VPWR VGND sg13g2_buf_8
Xfanout779 net781 net779 VPWR VGND sg13g2_buf_8
XFILLER_39_660 VPWR VGND sg13g2_fill_1
XFILLER_38_170 VPWR VGND sg13g2_fill_1
X_5009_ net159 VGND VPWR _0556_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\]
+ _0204_ sg13g2_dfrbpq_1
XFILLER_41_302 VPWR VGND sg13g2_decap_8
XFILLER_14_516 VPWR VGND sg13g2_fill_2
XFILLER_26_376 VPWR VGND sg13g2_fill_2
XFILLER_41_357 VPWR VGND sg13g2_fill_1
XFILLER_10_733 VPWR VGND sg13g2_fill_1
XFILLER_2_965 VPWR VGND sg13g2_decap_8
XFILLER_1_453 VPWR VGND sg13g2_fill_2
XFILLER_39_50 VPWR VGND sg13g2_fill_1
XFILLER_7_1003 VPWR VGND sg13g2_decap_8
XFILLER_39_72 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_fill_1
XFILLER_44_173 VPWR VGND sg13g2_fill_1
XFILLER_32_346 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_fill_2
XFILLER_9_553 VPWR VGND sg13g2_decap_8
X_2710_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\] _0741_ _0530_
+ VPWR VGND sg13g2_mux2_1
X_3690_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\] net583 _1420_ VPWR
+ VGND sg13g2_nor2_1
X_2641_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\] net789 _0724_ _0582_
+ VPWR VGND sg13g2_mux2_1
X_2572_ _0687_ _0682_ _0686_ VPWR VGND sg13g2_nand2_2
XFILLER_5_781 VPWR VGND sg13g2_fill_1
XFILLER_5_770 VPWR VGND sg13g2_decap_8
X_4311_ _2005_ _2009_ _2011_ VPWR VGND sg13g2_nor2_1
XFILLER_45_1020 VPWR VGND sg13g2_decap_4
X_4242_ _1948_ VPWR _1949_ VGND _0890_ _1945_ sg13g2_o21ai_1
X_4173_ _1786_ _1778_ _1896_ VPWR VGND sg13g2_xor2_1
X_3124_ _0799_ _0898_ _0904_ _0308_ VPWR VGND sg13g2_nor3_1
X_3055_ _0846_ tmds_green.dc_balancing_reg\[4\] net603 VPWR VGND sg13g2_nand2b_1
XFILLER_27_129 VPWR VGND sg13g2_decap_8
XFILLER_24_803 VPWR VGND sg13g2_decap_4
XFILLER_35_173 VPWR VGND sg13g2_fill_2
XFILLER_24_869 VPWR VGND sg13g2_decap_8
X_3957_ _1681_ _1680_ _1677_ _1683_ VPWR VGND sg13g2_a21o_1
XFILLER_23_368 VPWR VGND sg13g2_decap_4
Xclkbuf_0_clk_regs clk_regs clknet_0_clk_regs VPWR VGND sg13g2_buf_8
X_2908_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\] _0786_ _0294_
+ VPWR VGND sg13g2_mux2_1
X_3888_ _1617_ _1616_ _1449_ VPWR VGND sg13g2_nand2b_1
X_2839_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\] net783 _0770_ _0421_
+ VPWR VGND sg13g2_mux2_1
XFILLER_3_707 VPWR VGND sg13g2_fill_1
X_4509_ net675 net725 _0062_ VPWR VGND sg13g2_nor2_1
XFILLER_47_906 VPWR VGND sg13g2_decap_8
Xfanout565 net566 net565 VPWR VGND sg13g2_buf_8
Xfanout543 _0673_ net543 VPWR VGND sg13g2_buf_8
Xfanout554 net557 net554 VPWR VGND sg13g2_buf_8
XFILLER_46_405 VPWR VGND sg13g2_decap_4
Xfanout576 _0690_ net576 VPWR VGND sg13g2_buf_8
Xfanout587 net590 net587 VPWR VGND sg13g2_buf_8
Xfanout598 net599 net598 VPWR VGND sg13g2_buf_1
XFILLER_42_600 VPWR VGND sg13g2_decap_4
XFILLER_14_324 VPWR VGND sg13g2_decap_4
XFILLER_25_63 VPWR VGND sg13g2_decap_8
XFILLER_41_51 VPWR VGND sg13g2_decap_4
XFILLER_2_751 VPWR VGND sg13g2_decap_8
XFILLER_49_265 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_fill_1
XFILLER_18_630 VPWR VGND sg13g2_decap_4
XFILLER_18_663 VPWR VGND sg13g2_decap_8
XFILLER_17_173 VPWR VGND sg13g2_decap_8
XFILLER_18_685 VPWR VGND sg13g2_fill_2
XFILLER_18_696 VPWR VGND sg13g2_fill_1
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
X_4860_ net278 VGND VPWR _0411_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\]
+ _0068_ sg13g2_dfrbpq_1
XFILLER_20_305 VPWR VGND sg13g2_fill_1
X_3811_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\] net589 _1541_ VPWR
+ VGND sg13g2_nor2_1
X_4791_ net392 VGND VPWR _0342_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\]
+ _0042_ sg13g2_dfrbpq_1
XFILLER_20_316 VPWR VGND sg13g2_decap_8
XFILLER_20_338 VPWR VGND sg13g2_decap_8
X_3742_ _1471_ VPWR _1472_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\]
+ net585 sg13g2_o21ai_1
XFILLER_9_361 VPWR VGND sg13g2_decap_8
X_3673_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\] net554 _1403_ VPWR
+ VGND sg13g2_nor2_1
X_4872__251 VPWR VGND net251 sg13g2_tiehi
X_2624_ _0719_ _0713_ _0717_ VPWR VGND sg13g2_nand2_2
X_2555_ _0670_ _0667_ _0668_ _0669_ VPWR VGND sg13g2_and3_2
X_4225_ _1932_ tmds_red.dc_balancing_reg\[2\] _0883_ VPWR VGND sg13g2_xnor2_1
X_4156_ _1879_ _1877_ _1878_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_939 VPWR VGND sg13g2_decap_8
X_3107_ net569 _0894_ _0276_ VPWR VGND sg13g2_nor2_1
X_4087_ _1123_ _1807_ _1117_ _1810_ VPWR VGND sg13g2_nand3_1
XFILLER_37_983 VPWR VGND sg13g2_decap_8
X_3038_ _0808_ _0835_ _0001_ VPWR VGND sg13g2_nor2_1
XFILLER_36_460 VPWR VGND sg13g2_fill_1
XFILLER_12_828 VPWR VGND sg13g2_fill_2
X_4989_ net238 VGND VPWR _0536_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\]
+ _0184_ sg13g2_dfrbpq_1
XFILLER_20_883 VPWR VGND sg13g2_decap_8
XFILLER_3_537 VPWR VGND sg13g2_decap_4
XFILLER_11_98 VPWR VGND sg13g2_decap_4
XFILLER_4_1006 VPWR VGND sg13g2_decap_8
XFILLER_47_725 VPWR VGND sg13g2_fill_1
XFILLER_46_213 VPWR VGND sg13g2_decap_4
XFILLER_34_419 VPWR VGND sg13g2_fill_2
XFILLER_43_942 VPWR VGND sg13g2_decap_8
XFILLER_14_110 VPWR VGND sg13g2_fill_1
XFILLER_42_463 VPWR VGND sg13g2_fill_1
XFILLER_42_452 VPWR VGND sg13g2_decap_4
XFILLER_14_132 VPWR VGND sg13g2_fill_1
XFILLER_15_655 VPWR VGND sg13g2_fill_1
XFILLER_15_677 VPWR VGND sg13g2_decap_8
XFILLER_42_485 VPWR VGND sg13g2_fill_1
XFILLER_42_474 VPWR VGND sg13g2_fill_1
XFILLER_10_393 VPWR VGND sg13g2_fill_2
XFILLER_7_898 VPWR VGND sg13g2_decap_8
X_4010_ _1733_ _1732_ _1731_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_769 VPWR VGND sg13g2_fill_2
X_4912_ net172 VGND VPWR _0463_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\]
+ _0120_ sg13g2_dfrbpq_1
XFILLER_33_430 VPWR VGND sg13g2_decap_4
XFILLER_34_986 VPWR VGND sg13g2_decap_8
X_4843_ net311 VGND VPWR _0394_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\]
+ _0051_ sg13g2_dfrbpq_1
XFILLER_33_496 VPWR VGND sg13g2_fill_1
X_4774_ net54 VGND VPWR _0325_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\]
+ net633 sg13g2_dfrbpq_1
X_3725_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\] net588 _1455_ VPWR
+ VGND sg13g2_nor2_1
X_3656_ net592 _1380_ _1385_ _1386_ VPWR VGND sg13g2_nor3_1
X_2607_ net619 _0693_ _0709_ _0710_ VPWR VGND sg13g2_nor3_2
X_3587_ _1313_ _1314_ _1315_ _1316_ _1317_ VPWR VGND sg13g2_nor4_1
X_2538_ VPWR _0655_ net417 VGND sg13g2_inv_1
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_0_529 VPWR VGND sg13g2_fill_1
X_4811__352 VPWR VGND net352 sg13g2_tiehi
X_4208_ _0647_ net548 _1923_ VPWR VGND sg13g2_nor2_1
X_4139_ _1861_ VPWR _1862_ VGND _1840_ _1854_ sg13g2_o21ai_1
XFILLER_28_224 VPWR VGND sg13g2_fill_2
XFILLER_25_920 VPWR VGND sg13g2_decap_8
XFILLER_11_102 VPWR VGND sg13g2_fill_2
XFILLER_11_113 VPWR VGND sg13g2_decap_8
XFILLER_24_485 VPWR VGND sg13g2_decap_8
XFILLER_25_997 VPWR VGND sg13g2_decap_8
XFILLER_8_629 VPWR VGND sg13g2_fill_1
XFILLER_11_157 VPWR VGND sg13g2_fill_2
XFILLER_3_334 VPWR VGND sg13g2_fill_2
XFILLER_19_246 VPWR VGND sg13g2_decap_8
XFILLER_47_599 VPWR VGND sg13g2_fill_1
XFILLER_16_964 VPWR VGND sg13g2_decap_8
XFILLER_43_794 VPWR VGND sg13g2_fill_1
XFILLER_43_783 VPWR VGND sg13g2_fill_1
XFILLER_31_934 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_4
XFILLER_8_66 VPWR VGND sg13g2_decap_8
XFILLER_7_651 VPWR VGND sg13g2_decap_8
X_3510_ VPWR VGND _1227_ _1239_ _1237_ _1235_ _1240_ _1236_ sg13g2_a221oi_1
X_4490_ net652 net703 _0043_ VPWR VGND sg13g2_nor2_1
X_4793__388 VPWR VGND net388 sg13g2_tiehi
X_3441_ _1166_ _1168_ net545 _1171_ VPWR VGND sg13g2_nand3_1
X_3372_ _1102_ videogen.fancy_shader.n646\[7\] net629 VPWR VGND sg13g2_xnor2_1
X_5111_ net796 VGND VPWR serialize.n429\[8\] serialize.n417\[6\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_890 VPWR VGND sg13g2_decap_8
XFILLER_38_500 VPWR VGND sg13g2_decap_8
X_5042_ net205 VGND VPWR _0589_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\]
+ _0237_ sg13g2_dfrbpq_1
XFILLER_26_728 VPWR VGND sg13g2_fill_2
X_4908__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_22_956 VPWR VGND sg13g2_decap_8
X_4826_ net333 VGND VPWR _0377_ tmds_green.n126 net640 sg13g2_dfrbpq_2
X_4757_ net82 VGND VPWR _0308_ videogen.fancy_shader.video_x\[5\] net638 sg13g2_dfrbpq_2
X_3708_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\] net553 _1438_ VPWR
+ VGND sg13g2_nor2_1
X_4688_ net685 net735 _0241_ VPWR VGND sg13g2_nor2_1
X_3639_ net596 VPWR _1369_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\]
+ net562 sg13g2_o21ai_1
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_29_555 VPWR VGND sg13g2_decap_4
XFILLER_17_53 VPWR VGND sg13g2_decap_8
XFILLER_17_64 VPWR VGND sg13g2_fill_2
XFILLER_16_249 VPWR VGND sg13g2_decap_4
XFILLER_17_97 VPWR VGND sg13g2_fill_1
XFILLER_25_750 VPWR VGND sg13g2_fill_1
X_4922__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_13_923 VPWR VGND sg13g2_decap_8
XFILLER_40_775 VPWR VGND sg13g2_decap_4
XFILLER_8_415 VPWR VGND sg13g2_decap_8
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_decap_4
XFILLER_12_477 VPWR VGND sg13g2_fill_1
XFILLER_32_1011 VPWR VGND sg13g2_decap_8
XFILLER_8_459 VPWR VGND sg13g2_decap_4
X_4968__347 VPWR VGND net347 sg13g2_tiehi
X_5064__217 VPWR VGND net217 sg13g2_tiehi
Xhold4 serialize.n420\[0\] VPWR VGND net409 sg13g2_dlygate4sd3_1
XFILLER_47_352 VPWR VGND sg13g2_fill_2
XFILLER_47_341 VPWR VGND sg13g2_fill_2
XFILLER_35_514 VPWR VGND sg13g2_fill_1
X_3990_ _1716_ _1251_ _1715_ VPWR VGND sg13g2_nand2_1
X_2941_ videogen.fancy_shader.video_x\[5\] _0798_ _0799_ VPWR VGND sg13g2_and2_1
XFILLER_15_282 VPWR VGND sg13g2_decap_4
X_4611_ net691 net743 _0164_ VPWR VGND sg13g2_nor2_1
X_2872_ _0725_ _0772_ _0779_ VPWR VGND sg13g2_nor2_2
XFILLER_31_764 VPWR VGND sg13g2_fill_1
XFILLER_8_982 VPWR VGND sg13g2_decap_8
X_4542_ net679 net730 _0095_ VPWR VGND sg13g2_nor2_1
XFILLER_7_470 VPWR VGND sg13g2_decap_4
X_4473_ net661 net712 _0026_ VPWR VGND sg13g2_nor2_1
X_3424_ VGND VPWR _1136_ _1144_ _1154_ _1140_ sg13g2_a21oi_1
X_3355_ _1085_ _1084_ _1076_ VPWR VGND sg13g2_nand2b_1
X_3286_ _1016_ videogen.fancy_shader.n646\[2\] videogen.fancy_shader.video_x\[2\]
+ VPWR VGND sg13g2_xnor2_1
X_5025_ net365 VGND VPWR _0572_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\]
+ _0220_ sg13g2_dfrbpq_1
XFILLER_39_875 VPWR VGND sg13g2_decap_4
XFILLER_26_536 VPWR VGND sg13g2_fill_2
XFILLER_16_1006 VPWR VGND sg13g2_decap_8
XFILLER_10_926 VPWR VGND sg13g2_decap_8
XFILLER_22_775 VPWR VGND sg13g2_fill_2
X_4809_ net356 VGND VPWR _0360_ videogen.fancy_shader.video_y\[4\] net636 sg13g2_dfrbpq_2
XFILLER_0_123 VPWR VGND sg13g2_fill_1
XFILLER_0_156 VPWR VGND sg13g2_decap_8
XFILLER_45_867 VPWR VGND sg13g2_decap_4
XFILLER_44_333 VPWR VGND sg13g2_decap_8
XFILLER_17_558 VPWR VGND sg13g2_decap_8
XFILLER_13_720 VPWR VGND sg13g2_decap_8
XFILLER_32_528 VPWR VGND sg13g2_decap_8
XFILLER_32_539 VPWR VGND sg13g2_fill_2
XFILLER_40_594 VPWR VGND sg13g2_fill_1
XFILLER_12_285 VPWR VGND sg13g2_decap_8
XFILLER_8_267 VPWR VGND sg13g2_decap_8
XFILLER_8_289 VPWR VGND sg13g2_fill_1
XFILLER_5_974 VPWR VGND sg13g2_decap_8
XFILLER_5_56 VPWR VGND sg13g2_decap_8
X_4714__153 VPWR VGND net153 sg13g2_tiehi
X_3140_ _0914_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] _0915_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_39_138 VPWR VGND sg13g2_fill_2
X_3071_ _0861_ net548 _0860_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
X_3973_ _1699_ _1686_ _1698_ VPWR VGND sg13g2_nand2_1
X_2924_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\] net763 _0789_ _0281_
+ VPWR VGND sg13g2_mux2_1
X_2855_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\] _0775_ _0410_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_583 VPWR VGND sg13g2_fill_1
X_4525_ net658 net709 _0078_ VPWR VGND sg13g2_nor2_1
X_2786_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\] net788 _0757_ _0461_
+ VPWR VGND sg13g2_mux2_1
X_4456_ net569 _0894_ _0277_ VPWR VGND sg13g2_nor2_1
X_4387_ net604 _2001_ _2077_ _2078_ VPWR VGND sg13g2_nor3_1
X_3407_ _1067_ _1114_ _1132_ _1137_ VPWR VGND sg13g2_nor3_1
Xfanout703 net707 net703 VPWR VGND sg13g2_buf_8
Xfanout714 net724 net714 VPWR VGND sg13g2_buf_8
Xfanout725 net727 net725 VPWR VGND sg13g2_buf_8
X_3338_ _1068_ _1044_ _1058_ VPWR VGND sg13g2_nand2_1
Xfanout747 net749 net747 VPWR VGND sg13g2_buf_8
Xfanout736 net739 net736 VPWR VGND sg13g2_buf_1
Xfanout758 net759 net758 VPWR VGND sg13g2_buf_8
Xfanout769 net770 net769 VPWR VGND sg13g2_buf_8
X_3269_ videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\] videogen.fancy_shader.video_x\[7\]
+ _1000_ VPWR VGND _0902_ sg13g2_nand4_1
X_5008_ net163 VGND VPWR _0555_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\]
+ _0203_ sg13g2_dfrbpq_1
XFILLER_14_539 VPWR VGND sg13g2_decap_8
XFILLER_10_701 VPWR VGND sg13g2_decap_4
XFILLER_14_54 VPWR VGND sg13g2_fill_1
XFILLER_22_583 VPWR VGND sg13g2_decap_4
XFILLER_10_756 VPWR VGND sg13g2_decap_4
XFILLER_5_237 VPWR VGND sg13g2_fill_2
XFILLER_30_31 VPWR VGND sg13g2_fill_1
XFILLER_2_944 VPWR VGND sg13g2_decap_8
XFILLER_39_40 VPWR VGND sg13g2_fill_2
XFILLER_49_469 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_4
XFILLER_17_344 VPWR VGND sg13g2_fill_2
XFILLER_44_196 VPWR VGND sg13g2_fill_1
XFILLER_33_859 VPWR VGND sg13g2_decap_4
X_2640_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\] net775 _0724_ _0583_
+ VPWR VGND sg13g2_mux2_1
X_2571_ VGND VPWR _0685_ _0686_ _0672_ net600 sg13g2_a21oi_2
XFILLER_5_760 VPWR VGND sg13g2_fill_1
X_4310_ _2010_ _2009_ _2006_ VPWR VGND sg13g2_nand2b_1
XFILLER_4_292 VPWR VGND sg13g2_decap_8
X_4241_ _0891_ _1943_ _1944_ _1947_ _1948_ VPWR VGND sg13g2_or4_1
X_4172_ _1895_ _1177_ _1234_ VPWR VGND sg13g2_nand2_1
X_3123_ videogen.fancy_shader.video_x\[5\] _0798_ _0904_ VPWR VGND sg13g2_nor2_1
XFILLER_49_981 VPWR VGND sg13g2_decap_8
X_3054_ _0842_ net601 _0840_ _0845_ VPWR VGND sg13g2_mux2_1
XFILLER_36_620 VPWR VGND sg13g2_decap_4
XFILLER_35_130 VPWR VGND sg13g2_fill_1
XFILLER_36_642 VPWR VGND sg13g2_fill_2
XFILLER_36_653 VPWR VGND sg13g2_decap_4
XFILLER_35_141 VPWR VGND sg13g2_decap_4
XFILLER_36_686 VPWR VGND sg13g2_fill_2
X_3956_ _1680_ _1681_ _1682_ VPWR VGND sg13g2_and2_1
X_2907_ _0786_ _0688_ _0715_ VPWR VGND sg13g2_nand2_2
X_3887_ _1581_ VPWR _1616_ VGND _1599_ _1615_ sg13g2_o21ai_1
X_2838_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\] net773 _0770_ _0422_
+ VPWR VGND sg13g2_mux2_1
X_2769_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\] _0754_ _0475_
+ VPWR VGND sg13g2_mux2_1
X_4508_ net655 net706 _0061_ VPWR VGND sg13g2_nor2_1
X_4439_ tmds_blue.n193 _2077_ net604 _2128_ VPWR VGND sg13g2_nand3_1
Xfanout566 net567 net566 VPWR VGND sg13g2_buf_8
Xfanout544 _1055_ net544 VPWR VGND sg13g2_buf_8
Xfanout555 net557 net555 VPWR VGND sg13g2_buf_8
Xfanout588 net589 net588 VPWR VGND sg13g2_buf_8
Xfanout577 net578 net577 VPWR VGND sg13g2_buf_8
Xfanout599 _0638_ net599 VPWR VGND sg13g2_buf_8
XFILLER_46_439 VPWR VGND sg13g2_decap_4
X_5060__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_25_20 VPWR VGND sg13g2_fill_2
XFILLER_27_675 VPWR VGND sg13g2_decap_4
XFILLER_41_155 VPWR VGND sg13g2_decap_4
XFILLER_30_829 VPWR VGND sg13g2_fill_1
XFILLER_41_177 VPWR VGND sg13g2_decap_4
XFILLER_23_892 VPWR VGND sg13g2_decap_8
XFILLER_6_579 VPWR VGND sg13g2_decap_8
XFILLER_29_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_130 VPWR VGND sg13g2_decap_4
XFILLER_18_642 VPWR VGND sg13g2_fill_1
XFILLER_46_984 VPWR VGND sg13g2_decap_8
X_3810_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\] net580 _1540_ VPWR
+ VGND sg13g2_nor2_1
X_4790_ net394 VGND VPWR _0341_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\]
+ _0041_ sg13g2_dfrbpq_1
X_3741_ _1469_ _1470_ _1471_ VPWR VGND sg13g2_nor2_1
XFILLER_32_199 VPWR VGND sg13g2_fill_1
X_5037__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_9_340 VPWR VGND sg13g2_fill_2
XFILLER_13_391 VPWR VGND sg13g2_decap_8
X_5072__146 VPWR VGND net146 sg13g2_tiehi
X_3672_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\] net578 _1402_ VPWR
+ VGND sg13g2_nor2_1
X_2623_ VGND VPWR _0718_ _0701_ net577 sg13g2_or2_1
X_2554_ videogen.fancy_shader.video_x\[3\] videogen.fancy_shader.video_x\[2\] videogen.fancy_shader.video_x\[1\]
+ net630 _0669_ VPWR VGND sg13g2_nor4_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_5_590 VPWR VGND sg13g2_fill_2
X_4224_ VGND VPWR _0893_ _1930_ _0502_ _1931_ sg13g2_a21oi_1
X_4155_ _1858_ VPWR _1878_ VGND _1865_ _1868_ sg13g2_o21ai_1
XFILLER_29_918 VPWR VGND sg13g2_decap_8
XFILLER_28_417 VPWR VGND sg13g2_decap_8
X_3106_ _0894_ _0860_ _0893_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_951 VPWR VGND sg13g2_fill_2
X_4086_ _1808_ _1737_ _1809_ VPWR VGND sg13g2_xor2_1
X_3037_ _0835_ net794 _0807_ VPWR VGND sg13g2_nand2_1
XFILLER_23_133 VPWR VGND sg13g2_decap_8
XFILLER_24_667 VPWR VGND sg13g2_decap_8
XFILLER_23_177 VPWR VGND sg13g2_fill_1
X_4988_ net242 VGND VPWR _0535_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\]
+ _0183_ sg13g2_dfrbpq_1
X_3939_ _1665_ _1663_ _1664_ VPWR VGND sg13g2_nand2_1
X_5055__377 VPWR VGND net377 sg13g2_tiehi
X_4918__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_3_516 VPWR VGND sg13g2_decap_8
XFILLER_11_66 VPWR VGND sg13g2_fill_1
XFILLER_11_77 VPWR VGND sg13g2_decap_8
X_4734__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_19_406 VPWR VGND sg13g2_fill_2
XFILLER_19_439 VPWR VGND sg13g2_decap_4
XFILLER_43_921 VPWR VGND sg13g2_decap_8
XFILLER_27_450 VPWR VGND sg13g2_fill_1
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_fill_2
XFILLER_43_998 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_fill_2
X_4937__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_7_866 VPWR VGND sg13g2_decap_4
XFILLER_10_372 VPWR VGND sg13g2_fill_1
XFILLER_42_7 VPWR VGND sg13g2_decap_4
XFILLER_2_582 VPWR VGND sg13g2_fill_2
XFILLER_19_984 VPWR VGND sg13g2_decap_8
X_4911_ net174 VGND VPWR _0462_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\]
+ _0119_ sg13g2_dfrbpq_1
XFILLER_34_921 VPWR VGND sg13g2_decap_8
XFILLER_34_954 VPWR VGND sg13g2_fill_2
X_4842_ net313 VGND VPWR _0393_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\]
+ _0050_ sg13g2_dfrbpq_1
XFILLER_33_475 VPWR VGND sg13g2_decap_8
XFILLER_33_486 VPWR VGND sg13g2_fill_2
X_4773_ net56 VGND VPWR _0324_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[0\]
+ net633 sg13g2_dfrbpq_1
XFILLER_20_136 VPWR VGND sg13g2_decap_4
X_3724_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\] net579 _1454_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_181 VPWR VGND sg13g2_fill_2
X_3655_ _1381_ _1382_ _1383_ _1384_ _1385_ VPWR VGND sg13g2_nor4_1
X_2606_ net600 net543 net626 _0709_ VPWR VGND sg13g2_nand3_1
X_4954__393 VPWR VGND net393 sg13g2_tiehi
X_3586_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\] net551 _1316_ VPWR
+ VGND sg13g2_nor2_1
X_4207_ _0648_ _1922_ _0386_ VPWR VGND sg13g2_nor2_1
XFILLER_29_737 VPWR VGND sg13g2_decap_4
X_4138_ _1861_ _1830_ _1838_ VPWR VGND sg13g2_xnor2_1
X_4069_ VGND VPWR _1779_ _1785_ _1792_ _1786_ sg13g2_a21oi_1
X_4961__375 VPWR VGND net375 sg13g2_tiehi
XFILLER_24_453 VPWR VGND sg13g2_decap_4
XFILLER_25_976 VPWR VGND sg13g2_decap_8
XFILLER_4_825 VPWR VGND sg13g2_decap_4
XFILLER_19_225 VPWR VGND sg13g2_fill_1
XFILLER_47_578 VPWR VGND sg13g2_decap_8
XFILLER_16_943 VPWR VGND sg13g2_decap_8
XFILLER_15_442 VPWR VGND sg13g2_decap_8
XFILLER_31_913 VPWR VGND sg13g2_decap_8
XFILLER_8_89 VPWR VGND sg13g2_fill_1
XFILLER_11_681 VPWR VGND sg13g2_fill_1
XFILLER_11_692 VPWR VGND sg13g2_fill_2
XFILLER_7_696 VPWR VGND sg13g2_fill_2
XFILLER_6_195 VPWR VGND sg13g2_decap_4
X_3440_ _1165_ _1169_ _1170_ VPWR VGND sg13g2_nor2_1
XFILLER_40_4 VPWR VGND sg13g2_fill_1
X_3371_ videogen.fancy_shader.n646\[7\] net629 _1101_ VPWR VGND sg13g2_nor2_1
X_5110_ net796 VGND VPWR serialize.n429\[7\] serialize.n417\[5\] clknet_3_0__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5041_ net213 VGND VPWR _0588_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\]
+ _0236_ sg13g2_dfrbpq_1
XFILLER_26_2 VPWR VGND sg13g2_fill_1
XFILLER_38_578 VPWR VGND sg13g2_fill_2
XFILLER_22_935 VPWR VGND sg13g2_decap_8
XFILLER_34_795 VPWR VGND sg13g2_fill_2
X_4825_ net334 VGND VPWR _0376_ tmds_green.n100 net642 sg13g2_dfrbpq_2
XFILLER_21_456 VPWR VGND sg13g2_decap_4
XFILLER_21_478 VPWR VGND sg13g2_fill_1
X_4756_ net83 VGND VPWR _0307_ videogen.fancy_shader.video_x\[4\] net638 sg13g2_dfrbpq_2
X_4687_ net687 net738 _0240_ VPWR VGND sg13g2_nor2_1
X_3707_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\] net586 _1437_ VPWR
+ VGND sg13g2_nor2_1
X_3638_ _1364_ _1365_ _1366_ _1367_ _1368_ VPWR VGND sg13g2_nor4_1
X_3569_ net613 _1287_ _1298_ _1299_ VPWR VGND sg13g2_nor3_1
XFILLER_1_839 VPWR VGND sg13g2_decap_8
XFILLER_44_559 VPWR VGND sg13g2_decap_8
XFILLER_40_732 VPWR VGND sg13g2_decap_4
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_13_979 VPWR VGND sg13g2_decap_8
XFILLER_8_438 VPWR VGND sg13g2_fill_1
XFILLER_12_489 VPWR VGND sg13g2_decap_4
XFILLER_4_644 VPWR VGND sg13g2_fill_2
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_4_699 VPWR VGND sg13g2_fill_2
XFILLER_3_176 VPWR VGND sg13g2_fill_1
Xhold5 serialize.n420\[2\] VPWR VGND net410 sg13g2_dlygate4sd3_1
XFILLER_35_526 VPWR VGND sg13g2_decap_8
XFILLER_16_751 VPWR VGND sg13g2_decap_8
X_2940_ videogen.fancy_shader.video_x\[4\] _0796_ _0798_ VPWR VGND sg13g2_and2_1
X_2871_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[0\] net782 _0778_ _0397_
+ VPWR VGND sg13g2_mux2_1
X_4610_ net690 net744 _0163_ VPWR VGND sg13g2_nor2_1
XFILLER_30_286 VPWR VGND sg13g2_fill_1
XFILLER_8_961 VPWR VGND sg13g2_decap_8
X_4541_ net674 net726 _0094_ VPWR VGND sg13g2_nor2_1
X_4472_ net664 net715 _0025_ VPWR VGND sg13g2_nor2_1
X_3423_ _1151_ _1150_ _1148_ _1153_ VPWR VGND sg13g2_a21o_2
X_3354_ _1084_ _1080_ _1083_ VPWR VGND sg13g2_xnor2_1
X_3285_ _1015_ videogen.fancy_shader.n646\[2\] videogen.fancy_shader.video_x\[2\]
+ VPWR VGND sg13g2_nand2_1
X_5024_ net373 VGND VPWR _0571_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\]
+ _0219_ sg13g2_dfrbpq_1
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_38_320 VPWR VGND sg13g2_decap_8
XFILLER_0_1010 VPWR VGND sg13g2_decap_8
XFILLER_22_754 VPWR VGND sg13g2_decap_8
XFILLER_10_905 VPWR VGND sg13g2_decap_8
X_4808_ net358 VGND VPWR _0359_ videogen.fancy_shader.video_y\[3\] net636 sg13g2_dfrbpq_2
X_4739_ net113 VGND VPWR _0290_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\]
+ _0021_ sg13g2_dfrbpq_1
XFILLER_1_669 VPWR VGND sg13g2_decap_8
X_4852__294 VPWR VGND net294 sg13g2_tiehi
XFILLER_29_342 VPWR VGND sg13g2_fill_2
XFILLER_17_537 VPWR VGND sg13g2_fill_1
XFILLER_44_389 VPWR VGND sg13g2_decap_8
XFILLER_9_714 VPWR VGND sg13g2_decap_8
XFILLER_12_231 VPWR VGND sg13g2_decap_8
XFILLER_40_573 VPWR VGND sg13g2_fill_1
XFILLER_8_213 VPWR VGND sg13g2_fill_2
XFILLER_12_264 VPWR VGND sg13g2_fill_1
XFILLER_12_275 VPWR VGND sg13g2_fill_2
XFILLER_5_953 VPWR VGND sg13g2_decap_8
XFILLER_5_79 VPWR VGND sg13g2_fill_2
XFILLER_4_474 VPWR VGND sg13g2_fill_1
XFILLER_39_117 VPWR VGND sg13g2_decap_4
XFILLER_0_691 VPWR VGND sg13g2_decap_8
X_3070_ _0860_ tmds_red.n100 tmds_red.n102 VPWR VGND sg13g2_xnor2_1
XFILLER_36_813 VPWR VGND sg13g2_fill_1
XFILLER_39_1007 VPWR VGND sg13g2_decap_8
XFILLER_36_868 VPWR VGND sg13g2_fill_2
XFILLER_36_879 VPWR VGND sg13g2_decap_8
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_3972_ VGND VPWR _1695_ _1697_ _1698_ _1687_ sg13g2_a21oi_1
X_2923_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[3\] net752 _0789_ _0282_
+ VPWR VGND sg13g2_mux2_1
X_2854_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\] _0775_ _0411_
+ VPWR VGND sg13g2_mux2_1
X_2785_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\] net778 _0757_ _0462_
+ VPWR VGND sg13g2_mux2_1
X_4524_ net658 net708 _0077_ VPWR VGND sg13g2_nor2_1
X_4455_ _0642_ net569 _0272_ VPWR VGND sg13g2_nor2_1
Xfanout715 net718 net715 VPWR VGND sg13g2_buf_8
X_4386_ tmds_blue.n126 tmds_blue.n132 _2077_ VPWR VGND sg13g2_and2_1
X_3406_ VGND VPWR _1136_ _1135_ _1134_ sg13g2_or2_1
Xfanout704 net706 net704 VPWR VGND sg13g2_buf_8
Xfanout737 net738 net737 VPWR VGND sg13g2_buf_8
Xfanout726 net727 net726 VPWR VGND sg13g2_buf_8
X_3337_ VPWR _1067_ _1066_ VGND sg13g2_inv_1
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_1
Xfanout759 net760 net759 VPWR VGND sg13g2_buf_8
X_3268_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[3\] _0998_ _0369_ _0999_
+ sg13g2_a21oi_1
XFILLER_39_695 VPWR VGND sg13g2_decap_4
XFILLER_39_673 VPWR VGND sg13g2_decap_8
X_3199_ _0951_ _0955_ _0336_ VPWR VGND sg13g2_nor2_1
X_4882__232 VPWR VGND net232 sg13g2_tiehi
X_5007_ net167 VGND VPWR _0554_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\]
+ _0202_ sg13g2_dfrbpq_1
XFILLER_27_813 VPWR VGND sg13g2_decap_4
X_4808__358 VPWR VGND net358 sg13g2_tiehi
XFILLER_14_518 VPWR VGND sg13g2_fill_1
XFILLER_22_562 VPWR VGND sg13g2_decap_8
XFILLER_10_713 VPWR VGND sg13g2_decap_4
XFILLER_14_66 VPWR VGND sg13g2_decap_8
XFILLER_14_99 VPWR VGND sg13g2_decap_8
XFILLER_6_728 VPWR VGND sg13g2_fill_1
XFILLER_2_923 VPWR VGND sg13g2_decap_8
XFILLER_39_30 VPWR VGND sg13g2_decap_4
XFILLER_1_455 VPWR VGND sg13g2_fill_1
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_49_426 VPWR VGND sg13g2_decap_8
XFILLER_17_301 VPWR VGND sg13g2_fill_2
XFILLER_45_632 VPWR VGND sg13g2_decap_4
XFILLER_18_846 VPWR VGND sg13g2_decap_4
X_4744__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_32_359 VPWR VGND sg13g2_decap_8
XFILLER_40_370 VPWR VGND sg13g2_fill_2
XFILLER_13_573 VPWR VGND sg13g2_fill_1
X_2570_ VPWR _0685_ _0684_ VGND sg13g2_inv_1
XFILLER_5_794 VPWR VGND sg13g2_decap_8
X_4240_ _1929_ _1942_ _1947_ VPWR VGND sg13g2_and2_1
X_4171_ _1885_ _1886_ _1889_ _1893_ _1894_ VPWR VGND sg13g2_nor4_1
X_3122_ _0798_ _0903_ _0307_ VPWR VGND sg13g2_nor2_1
XFILLER_49_960 VPWR VGND sg13g2_decap_8
X_3053_ _0844_ net602 _0840_ VPWR VGND sg13g2_nand2_2
XFILLER_17_890 VPWR VGND sg13g2_decap_4
XFILLER_23_348 VPWR VGND sg13g2_decap_4
XFILLER_24_849 VPWR VGND sg13g2_decap_4
XFILLER_35_175 VPWR VGND sg13g2_fill_1
XFILLER_36_698 VPWR VGND sg13g2_decap_8
X_3955_ _1658_ _1672_ _1679_ _1681_ VPWR VGND sg13g2_or3_1
XFILLER_32_860 VPWR VGND sg13g2_decap_8
X_2906_ net785 videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\] _0785_ _0295_
+ VPWR VGND sg13g2_mux2_1
X_3886_ net2 VPWR _1615_ VGND videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\]
+ _1614_ sg13g2_o21ai_1
XFILLER_31_381 VPWR VGND sg13g2_decap_8
X_2837_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\] net763 _0770_ _0423_
+ VPWR VGND sg13g2_mux2_1
X_2768_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\] _0754_ _0476_
+ VPWR VGND sg13g2_mux2_1
X_2699_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\] _0739_ _0539_
+ VPWR VGND sg13g2_mux2_1
X_4507_ net668 net720 _0060_ VPWR VGND sg13g2_nor2_1
X_4438_ _2116_ VPWR _2127_ VGND _2115_ _2118_ sg13g2_o21ai_1
X_4369_ _2063_ _0847_ _2062_ VPWR VGND sg13g2_nand2_1
Xfanout545 _1021_ net545 VPWR VGND sg13g2_buf_8
Xfanout556 net557 net556 VPWR VGND sg13g2_buf_8
Xfanout589 net590 net589 VPWR VGND sg13g2_buf_8
Xfanout578 net581 net578 VPWR VGND sg13g2_buf_8
Xfanout567 net568 net567 VPWR VGND sg13g2_buf_8
XFILLER_27_654 VPWR VGND sg13g2_fill_2
XFILLER_26_131 VPWR VGND sg13g2_fill_2
XFILLER_15_849 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_26_175 VPWR VGND sg13g2_fill_2
XFILLER_41_134 VPWR VGND sg13g2_decap_8
XFILLER_14_348 VPWR VGND sg13g2_fill_2
XFILLER_14_359 VPWR VGND sg13g2_fill_1
XFILLER_23_871 VPWR VGND sg13g2_decap_8
XFILLER_10_521 VPWR VGND sg13g2_decap_4
XFILLER_6_525 VPWR VGND sg13g2_decap_8
XFILLER_6_558 VPWR VGND sg13g2_fill_1
XFILLER_2_775 VPWR VGND sg13g2_fill_2
XFILLER_1_274 VPWR VGND sg13g2_decap_8
XFILLER_38_919 VPWR VGND sg13g2_decap_8
XFILLER_49_289 VPWR VGND sg13g2_decap_8
XFILLER_46_963 VPWR VGND sg13g2_decap_8
XFILLER_17_142 VPWR VGND sg13g2_decap_8
XFILLER_17_153 VPWR VGND sg13g2_fill_1
XFILLER_18_687 VPWR VGND sg13g2_fill_1
XFILLER_33_602 VPWR VGND sg13g2_fill_1
XFILLER_45_495 VPWR VGND sg13g2_fill_2
XFILLER_45_484 VPWR VGND sg13g2_decap_8
X_3740_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\] net561 _1470_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_14_893 VPWR VGND sg13g2_fill_2
X_3671_ net597 VPWR _1401_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\]
+ net563 sg13g2_o21ai_1
X_2622_ net578 _0701_ _0717_ VPWR VGND sg13g2_nor2_2
X_2553_ videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\] videogen.fancy_shader.video_x\[4\]
+ _0668_ VPWR VGND sg13g2_nor3_1
X_4223_ _0836_ VPWR _1931_ VGND _0893_ _1930_ sg13g2_o21ai_1
X_4154_ _1877_ _1839_ _1854_ VPWR VGND sg13g2_xnor2_1
X_4085_ _1808_ _1117_ _1807_ VPWR VGND sg13g2_nand2_1
X_3105_ net570 _0893_ _0275_ VPWR VGND sg13g2_nor2_1
X_3036_ VPWR clk_video _0006_ VGND sg13g2_inv_1
XFILLER_36_451 VPWR VGND sg13g2_decap_4
XFILLER_23_112 VPWR VGND sg13g2_decap_8
XFILLER_24_613 VPWR VGND sg13g2_fill_1
XFILLER_24_646 VPWR VGND sg13g2_fill_1
X_4987_ net246 VGND VPWR _0534_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\]
+ _0182_ sg13g2_dfrbpq_1
X_3938_ _1664_ _1653_ _1655_ VPWR VGND sg13g2_nand2_1
X_3869_ VPWR VGND net597 net613 _1597_ _1593_ _1598_ _1596_ sg13g2_a221oi_1
XFILLER_46_237 VPWR VGND sg13g2_decap_8
X_4849__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_43_900 VPWR VGND sg13g2_decap_8
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_43_977 VPWR VGND sg13g2_decap_8
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_14_167 VPWR VGND sg13g2_decap_8
XFILLER_14_178 VPWR VGND sg13g2_fill_2
XFILLER_30_616 VPWR VGND sg13g2_decap_4
XFILLER_11_885 VPWR VGND sg13g2_fill_2
XFILLER_6_377 VPWR VGND sg13g2_fill_2
XFILLER_42_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_963 VPWR VGND sg13g2_decap_8
XFILLER_46_782 VPWR VGND sg13g2_decap_8
XFILLER_18_495 VPWR VGND sg13g2_decap_4
X_4910_ net176 VGND VPWR _0461_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\]
+ _0118_ sg13g2_dfrbpq_1
X_4841_ net315 VGND VPWR _0392_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\]
+ _0049_ sg13g2_dfrbpq_1
XFILLER_20_104 VPWR VGND sg13g2_decap_4
XFILLER_21_638 VPWR VGND sg13g2_decap_8
XFILLER_33_465 VPWR VGND sg13g2_decap_4
X_4772_ net58 VGND VPWR _0323_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ net631 sg13g2_dfrbpq_1
X_3723_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\] net555 _1453_ VPWR
+ VGND sg13g2_nor2_1
X_3654_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\] net550 _1384_ VPWR
+ VGND sg13g2_nor2_1
X_2605_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\] _0708_ _0602_
+ VPWR VGND sg13g2_mux2_1
X_3585_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\] net575 _1315_ VPWR
+ VGND sg13g2_nor2_1
X_2536_ VPWR _0654_ tmds_red.dc_balancing_reg\[2\] VGND sg13g2_inv_1
X_4206_ VGND VPWR _0884_ _1917_ _1922_ _1921_ sg13g2_a21oi_1
XFILLER_3_90 VPWR VGND sg13g2_decap_8
X_4137_ _1860_ _1854_ _1855_ _1859_ VPWR VGND sg13g2_and3_1
X_4068_ _1790_ _1789_ _1177_ _1791_ VPWR VGND sg13g2_a21o_1
X_3019_ net422 green_tmds_par\[2\] net697 serialize.n428\[4\] VPWR VGND sg13g2_mux2_1
XFILLER_19_1005 VPWR VGND sg13g2_decap_8
XFILLER_25_955 VPWR VGND sg13g2_decap_8
X_5018__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_36_292 VPWR VGND sg13g2_decap_4
X_4879__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_12_638 VPWR VGND sg13g2_fill_1
XFILLER_11_159 VPWR VGND sg13g2_fill_1
XFILLER_22_11 VPWR VGND sg13g2_decap_4
XFILLER_22_66 VPWR VGND sg13g2_fill_1
XFILLER_3_336 VPWR VGND sg13g2_fill_1
XFILLER_3_347 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_16_922 VPWR VGND sg13g2_decap_8
X_4862__274 VPWR VGND net274 sg13g2_tiehi
XFILLER_15_421 VPWR VGND sg13g2_decap_8
XFILLER_43_774 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_fill_2
XFILLER_16_999 VPWR VGND sg13g2_decap_8
XFILLER_8_24 VPWR VGND sg13g2_fill_1
X_4768__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_30_424 VPWR VGND sg13g2_fill_1
XFILLER_31_969 VPWR VGND sg13g2_decap_8
X_4783__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_8_79 VPWR VGND sg13g2_decap_4
XFILLER_10_181 VPWR VGND sg13g2_fill_2
XFILLER_6_174 VPWR VGND sg13g2_decap_8
X_3370_ _1100_ net610 videogen.fancy_shader.video_x\[8\] VPWR VGND sg13g2_nand2_1
X_5040_ net221 VGND VPWR _0587_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\]
+ _0235_ sg13g2_dfrbpq_1
XFILLER_46_590 VPWR VGND sg13g2_decap_4
XFILLER_34_752 VPWR VGND sg13g2_decap_4
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_21_435 VPWR VGND sg13g2_decap_8
X_4824_ net335 VGND VPWR _0375_ tmds_blue.n132 net640 sg13g2_dfrbpq_2
X_4755_ net84 VGND VPWR _0306_ videogen.fancy_shader.video_x\[3\] net637 sg13g2_dfrbpq_2
X_3706_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\] net565 _1436_ VPWR
+ VGND sg13g2_nor2_1
X_4686_ net685 net735 _0239_ VPWR VGND sg13g2_nor2_1
XFILLER_49_1009 VPWR VGND sg13g2_decap_8
X_3637_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\] net551 _1367_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_1_818 VPWR VGND sg13g2_decap_8
X_3568_ net618 _1292_ _1297_ _1298_ VPWR VGND sg13g2_nor3_1
X_2519_ _0637_ net612 VPWR VGND sg13g2_inv_2
X_3499_ _1217_ _1215_ _1229_ VPWR VGND sg13g2_xor2_1
XFILLER_29_579 VPWR VGND sg13g2_decap_8
XFILLER_44_516 VPWR VGND sg13g2_fill_1
XFILLER_17_66 VPWR VGND sg13g2_fill_1
XFILLER_17_88 VPWR VGND sg13g2_decap_8
XFILLER_24_240 VPWR VGND sg13g2_decap_4
XFILLER_25_785 VPWR VGND sg13g2_fill_1
XFILLER_13_958 VPWR VGND sg13g2_decap_8
XFILLER_33_54 VPWR VGND sg13g2_fill_1
XFILLER_33_65 VPWR VGND sg13g2_decap_8
XFILLER_33_76 VPWR VGND sg13g2_fill_2
X_4892__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_4_623 VPWR VGND sg13g2_fill_2
XFILLER_3_122 VPWR VGND sg13g2_decap_4
X_4792__390 VPWR VGND net390 sg13g2_tiehi
XFILLER_3_166 VPWR VGND sg13g2_decap_4
XFILLER_0_884 VPWR VGND sg13g2_decap_8
Xhold6 serialize.n420\[3\] VPWR VGND net411 sg13g2_dlygate4sd3_1
XFILLER_12_9 VPWR VGND sg13g2_decap_8
XFILLER_48_888 VPWR VGND sg13g2_decap_8
XFILLER_47_365 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_fill_1
XFILLER_47_387 VPWR VGND sg13g2_fill_2
XFILLER_28_590 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
X_2870_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[1\] net772 _0778_ _0398_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_796 VPWR VGND sg13g2_decap_4
XFILLER_8_940 VPWR VGND sg13g2_decap_8
X_4540_ net679 net730 _0093_ VPWR VGND sg13g2_nor2_1
X_5020__51 VPWR VGND net51 sg13g2_tiehi
X_4471_ net662 net713 _0024_ VPWR VGND sg13g2_nor2_1
X_3422_ _1152_ _1150_ _1151_ VPWR VGND sg13g2_nand2_1
X_3353_ _1083_ _1082_ _1081_ VPWR VGND sg13g2_nand2b_1
X_3284_ _1011_ VPWR _1014_ VGND _1012_ _1013_ sg13g2_o21ai_1
X_5023_ net381 VGND VPWR _0570_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\]
+ _0218_ sg13g2_dfrbpq_1
XFILLER_38_332 VPWR VGND sg13g2_decap_4
XFILLER_22_722 VPWR VGND sg13g2_decap_8
XFILLER_22_733 VPWR VGND sg13g2_fill_1
X_4807_ net360 VGND VPWR _0358_ videogen.fancy_shader.video_y\[2\] net636 sg13g2_dfrbpq_2
X_2999_ net700 net410 serialize.n431\[2\] VPWR VGND sg13g2_nor2b_1
X_4738_ net115 VGND VPWR _0289_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\]
+ _0020_ sg13g2_dfrbpq_1
X_4669_ net687 net738 _0222_ VPWR VGND sg13g2_nor2_1
X_5013__118 VPWR VGND net118 sg13g2_tiehi
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_43 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_fill_1
XFILLER_25_582 VPWR VGND sg13g2_decap_8
XFILLER_25_593 VPWR VGND sg13g2_fill_1
XFILLER_44_97 VPWR VGND sg13g2_decap_4
XFILLER_13_755 VPWR VGND sg13g2_decap_8
XFILLER_40_585 VPWR VGND sg13g2_fill_1
XFILLER_9_748 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_5_932 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_fill_1
X_5068__185 VPWR VGND net185 sg13g2_tiehi
X_4929__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_0_670 VPWR VGND sg13g2_decap_8
XFILLER_48_641 VPWR VGND sg13g2_decap_8
XFILLER_47_162 VPWR VGND sg13g2_fill_2
XFILLER_47_151 VPWR VGND sg13g2_fill_1
X_3971_ _1697_ _1683_ _1696_ VPWR VGND sg13g2_nand2_1
X_2922_ _0699_ _0772_ _0789_ VPWR VGND sg13g2_nor2_2
X_2853_ net756 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\] _0775_ _0412_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_574 VPWR VGND sg13g2_decap_8
X_2784_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\] net771 _0757_ _0463_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_781 VPWR VGND sg13g2_decap_8
X_4523_ net675 net709 _0076_ VPWR VGND sg13g2_nor2_1
X_4454_ net679 net730 _0009_ VPWR VGND sg13g2_nor2_1
X_3405_ _1135_ net544 _1127_ VPWR VGND sg13g2_nand2_1
Xfanout705 net706 net705 VPWR VGND sg13g2_buf_1
X_4385_ tmds_blue.n193 tmds_blue.n132 _2076_ VPWR VGND sg13g2_xor2_1
Xfanout716 net718 net716 VPWR VGND sg13g2_buf_1
X_3336_ _1064_ _1065_ _1066_ VPWR VGND sg13g2_and2_1
Xfanout727 net734 net727 VPWR VGND sg13g2_buf_2
Xfanout749 _0648_ net749 VPWR VGND sg13g2_buf_8
Xfanout738 net739 net738 VPWR VGND sg13g2_buf_8
X_5006_ net171 VGND VPWR _0553_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\]
+ _0201_ sg13g2_dfrbpq_1
XFILLER_22_1012 VPWR VGND sg13g2_decap_8
X_3267_ net793 VPWR _0999_ VGND videogen.test_lut_thingy.gol_counter_reg\[3\] _0998_
+ sg13g2_o21ai_1
X_3198_ _0955_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] _0954_ VPWR
+ VGND sg13g2_xnor2_1
XFILLER_38_195 VPWR VGND sg13g2_decap_4
XFILLER_26_346 VPWR VGND sg13g2_decap_8
XFILLER_41_316 VPWR VGND sg13g2_decap_4
XFILLER_14_89 VPWR VGND sg13g2_fill_2
XFILLER_5_239 VPWR VGND sg13g2_fill_1
XFILLER_2_902 VPWR VGND sg13g2_decap_8
XFILLER_7_1017 VPWR VGND sg13g2_decap_8
XFILLER_2_979 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_86 VPWR VGND sg13g2_fill_2
XFILLER_17_346 VPWR VGND sg13g2_fill_1
XFILLER_44_154 VPWR VGND sg13g2_fill_1
XFILLER_33_806 VPWR VGND sg13g2_decap_8
XFILLER_33_817 VPWR VGND sg13g2_fill_1
XFILLER_44_187 VPWR VGND sg13g2_decap_8
XFILLER_26_891 VPWR VGND sg13g2_decap_8
XFILLER_9_512 VPWR VGND sg13g2_decap_8
XFILLER_9_567 VPWR VGND sg13g2_fill_2
XFILLER_9_578 VPWR VGND sg13g2_fill_1
X_4170_ _1893_ _1890_ _1892_ VPWR VGND sg13g2_xnor2_1
X_3121_ _0903_ net795 _0902_ VPWR VGND sg13g2_nand2_1
XFILLER_48_471 VPWR VGND sg13g2_decap_4
X_3052_ _0843_ tmds_green.n100 _0642_ VPWR VGND sg13g2_nand2_1
XFILLER_48_493 VPWR VGND sg13g2_decap_8
XFILLER_35_121 VPWR VGND sg13g2_decap_8
XFILLER_24_828 VPWR VGND sg13g2_decap_8
XFILLER_23_327 VPWR VGND sg13g2_decap_8
XFILLER_35_198 VPWR VGND sg13g2_decap_4
X_3954_ _1679_ VPWR _1680_ VGND _1658_ _1672_ sg13g2_o21ai_1
X_2905_ net773 videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\] _0785_ _0296_
+ VPWR VGND sg13g2_mux2_1
X_3885_ _1613_ VPWR _1614_ VGND net612 _1604_ sg13g2_o21ai_1
X_2836_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\] net753 _0770_ _0424_
+ VPWR VGND sg13g2_mux2_1
X_2767_ _0754_ _0710_ _0720_ VPWR VGND sg13g2_nand2_2
X_2698_ net766 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\] _0739_ _0540_
+ VPWR VGND sg13g2_mux2_1
X_4506_ net659 net710 _0059_ VPWR VGND sg13g2_nor2_1
X_4437_ VGND VPWR _2121_ _2126_ _0626_ net571 sg13g2_a21oi_1
X_4368_ _2062_ _2050_ _2054_ VPWR VGND sg13g2_xnor2_1
Xfanout546 _1031_ net546 VPWR VGND sg13g2_buf_8
Xfanout557 net558 net557 VPWR VGND sg13g2_buf_8
X_4299_ _1998_ _2000_ _0612_ VPWR VGND sg13g2_nor2_1
Xfanout568 _1253_ net568 VPWR VGND sg13g2_buf_8
X_3319_ VPWR VGND _1047_ _1048_ _1007_ videogen.fancy_shader.video_y\[3\] _1049_ net611
+ sg13g2_a221oi_1
Xfanout579 net581 net579 VPWR VGND sg13g2_buf_8
X_4964__363 VPWR VGND net363 sg13g2_tiehi
XFILLER_27_600 VPWR VGND sg13g2_decap_8
XFILLER_27_622 VPWR VGND sg13g2_fill_2
XFILLER_14_338 VPWR VGND sg13g2_decap_4
XFILLER_26_187 VPWR VGND sg13g2_decap_8
XFILLER_26_198 VPWR VGND sg13g2_fill_1
X_4971__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_10_566 VPWR VGND sg13g2_fill_1
XFILLER_41_87 VPWR VGND sg13g2_fill_2
XFILLER_2_765 VPWR VGND sg13g2_fill_2
XFILLER_49_224 VPWR VGND sg13g2_decap_4
XFILLER_49_202 VPWR VGND sg13g2_decap_8
XFILLER_2_787 VPWR VGND sg13g2_decap_8
XFILLER_49_279 VPWR VGND sg13g2_decap_4
XFILLER_46_942 VPWR VGND sg13g2_decap_8
XFILLER_45_474 VPWR VGND sg13g2_decap_4
XFILLER_17_187 VPWR VGND sg13g2_fill_2
XFILLER_32_102 VPWR VGND sg13g2_decap_4
XFILLER_33_614 VPWR VGND sg13g2_decap_4
XFILLER_32_146 VPWR VGND sg13g2_fill_2
XFILLER_9_342 VPWR VGND sg13g2_fill_1
XFILLER_9_353 VPWR VGND sg13g2_decap_4
X_3670_ _1399_ VPWR _1400_ VGND _1363_ _1375_ sg13g2_o21ai_1
X_2621_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\] _0716_ _0594_
+ VPWR VGND sg13g2_mux2_1
X_2552_ net629 _0666_ _0667_ VPWR VGND sg13g2_and2_1
XFILLER_5_592 VPWR VGND sg13g2_fill_1
X_4222_ VPWR _1930_ _1929_ VGND sg13g2_inv_1
X_4153_ _1857_ _1870_ _1871_ _1875_ _1876_ VPWR VGND sg13g2_nor4_1
X_4084_ _1052_ _1063_ _1084_ _1799_ _1807_ VPWR VGND sg13g2_and4_1
X_3104_ _0890_ _0889_ net548 _0893_ VPWR VGND sg13g2_mux2_1
XFILLER_37_953 VPWR VGND sg13g2_fill_1
X_3035_ net679 net730 _0006_ VPWR VGND sg13g2_nor2_1
XFILLER_37_997 VPWR VGND sg13g2_decap_8
X_4986_ net250 VGND VPWR _0533_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\]
+ _0181_ sg13g2_dfrbpq_1
X_3937_ _1648_ VPWR _1663_ VGND _1652_ _1656_ sg13g2_o21ai_1
XFILLER_23_157 VPWR VGND sg13g2_fill_2
XFILLER_32_691 VPWR VGND sg13g2_fill_1
X_3868_ _1580_ VPWR _1597_ VGND _1571_ _1575_ sg13g2_o21ai_1
X_2819_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\] net788 _0766_ _0437_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_897 VPWR VGND sg13g2_fill_2
X_3799_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[3\] net586 _1529_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_19_408 VPWR VGND sg13g2_fill_1
XFILLER_19_419 VPWR VGND sg13g2_fill_2
XFILLER_28_942 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_36_32 VPWR VGND sg13g2_fill_2
XFILLER_43_956 VPWR VGND sg13g2_decap_8
XFILLER_6_334 VPWR VGND sg13g2_fill_2
XFILLER_38_717 VPWR VGND sg13g2_decap_4
XFILLER_19_942 VPWR VGND sg13g2_decap_8
XFILLER_46_761 VPWR VGND sg13g2_decap_4
XFILLER_34_945 VPWR VGND sg13g2_fill_1
X_4840_ net317 VGND VPWR _0391_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\]
+ _0048_ sg13g2_dfrbpq_1
XFILLER_34_956 VPWR VGND sg13g2_fill_1
X_4771_ net60 VGND VPWR _0322_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\]
+ net631 sg13g2_dfrbpq_1
X_3722_ net618 VPWR _1452_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\]
+ net565 sg13g2_o21ai_1
XFILLER_9_194 VPWR VGND sg13g2_decap_8
X_3653_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\] net573 _1383_ VPWR
+ VGND sg13g2_nor2_1
X_2604_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\] _0708_ _0603_
+ VPWR VGND sg13g2_mux2_1
X_3584_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\] net585 _1314_ VPWR
+ VGND sg13g2_nor2_1
X_2535_ VPWR _0653_ tmds_red.dc_balancing_reg\[3\] VGND sg13g2_inv_1
X_4205_ _1920_ VPWR _1921_ VGND _1916_ _1918_ sg13g2_o21ai_1
X_4136_ _1798_ _1840_ _1859_ VPWR VGND sg13g2_nor2_1
XFILLER_29_728 VPWR VGND sg13g2_fill_1
X_4067_ _1790_ _1234_ _1778_ VPWR VGND sg13g2_nand2_1
X_3018_ _0834_ VPWR serialize.n428\[3\] VGND _0656_ net697 sg13g2_o21ai_1
XFILLER_24_400 VPWR VGND sg13g2_fill_1
XFILLER_25_934 VPWR VGND sg13g2_decap_8
XFILLER_40_904 VPWR VGND sg13g2_fill_2
XFILLER_40_937 VPWR VGND sg13g2_decap_4
XFILLER_24_466 VPWR VGND sg13g2_decap_4
X_4969_ net320 VGND VPWR _0516_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\]
+ _0164_ sg13g2_dfrbpq_1
XFILLER_11_127 VPWR VGND sg13g2_decap_8
XFILLER_22_78 VPWR VGND sg13g2_decap_8
XFILLER_3_359 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_16_978 VPWR VGND sg13g2_decap_8
XFILLER_30_447 VPWR VGND sg13g2_decap_8
XFILLER_31_948 VPWR VGND sg13g2_decap_8
XFILLER_30_458 VPWR VGND sg13g2_fill_1
XFILLER_7_610 VPWR VGND sg13g2_fill_2
XFILLER_7_665 VPWR VGND sg13g2_fill_2
XFILLER_2_370 VPWR VGND sg13g2_decap_8
XFILLER_2_381 VPWR VGND sg13g2_fill_1
XFILLER_2_392 VPWR VGND sg13g2_decap_8
XFILLER_38_536 VPWR VGND sg13g2_decap_4
X_4841__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_34_731 VPWR VGND sg13g2_fill_1
XFILLER_21_403 VPWR VGND sg13g2_decap_8
XFILLER_33_263 VPWR VGND sg13g2_fill_1
XFILLER_34_764 VPWR VGND sg13g2_decap_4
X_4823_ net336 VGND VPWR _0374_ tmds_blue.n126 net640 sg13g2_dfrbpq_1
XFILLER_34_797 VPWR VGND sg13g2_fill_1
X_4754_ net85 VGND VPWR _0305_ videogen.fancy_shader.video_x\[2\] net637 sg13g2_dfrbpq_2
XFILLER_21_469 VPWR VGND sg13g2_decap_8
X_3705_ net618 VPWR _1435_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\]
+ net577 sg13g2_o21ai_1
X_4685_ net687 net739 _0238_ VPWR VGND sg13g2_nor2_1
X_3636_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\] net575 _1366_ VPWR
+ VGND sg13g2_nor2_1
X_3567_ _1293_ _1294_ _1295_ _1296_ _1297_ VPWR VGND sg13g2_nor4_1
X_2518_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _0636_ VPWR VGND sg13g2_inv_4
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_3498_ _1219_ _1227_ _1228_ VPWR VGND sg13g2_nor2_1
X_5099_ net800 VGND VPWR serialize.n431\[4\] serialize.n420\[2\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4119_ _1842_ _1771_ _1841_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_23 VPWR VGND sg13g2_fill_2
XFILLER_17_709 VPWR VGND sg13g2_decap_8
XFILLER_44_528 VPWR VGND sg13g2_decap_8
XFILLER_12_414 VPWR VGND sg13g2_decap_4
XFILLER_12_425 VPWR VGND sg13g2_fill_2
XFILLER_13_937 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_fill_2
XFILLER_33_22 VPWR VGND sg13g2_fill_1
XFILLER_8_429 VPWR VGND sg13g2_fill_2
XFILLER_21_992 VPWR VGND sg13g2_decap_8
XFILLER_4_646 VPWR VGND sg13g2_fill_1
X_4933__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_0_863 VPWR VGND sg13g2_decap_8
Xhold7 serialize.n420\[4\] VPWR VGND net412 sg13g2_dlygate4sd3_1
XFILLER_48_867 VPWR VGND sg13g2_decap_8
XFILLER_35_506 VPWR VGND sg13g2_fill_2
XFILLER_15_230 VPWR VGND sg13g2_fill_2
XFILLER_31_723 VPWR VGND sg13g2_fill_1
XFILLER_12_981 VPWR VGND sg13g2_decap_8
XFILLER_7_440 VPWR VGND sg13g2_fill_2
X_4470_ net664 net715 _0023_ VPWR VGND sg13g2_nor2_1
XFILLER_8_996 VPWR VGND sg13g2_decap_8
X_3421_ _1127_ VPWR _1151_ VGND _1133_ _1149_ sg13g2_o21ai_1
XFILLER_48_1021 VPWR VGND sg13g2_decap_8
X_3352_ VGND VPWR _1082_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.video_y\[6\]
+ sg13g2_or2_1
XFILLER_39_812 VPWR VGND sg13g2_fill_2
X_3283_ _1013_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_x\[1\]
+ VPWR VGND sg13g2_xnor2_1
X_5022_ net35 VGND VPWR _0569_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\]
+ _0217_ sg13g2_dfrbpq_1
XFILLER_17_0 VPWR VGND sg13g2_decap_4
X_4806_ net362 VGND VPWR _0357_ videogen.fancy_shader.video_y\[1\] net637 sg13g2_dfrbpq_2
X_2998_ net699 net408 serialize.n431\[1\] VPWR VGND sg13g2_nor2b_1
XFILLER_22_789 VPWR VGND sg13g2_decap_8
X_4737_ net117 VGND VPWR _0288_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\]
+ _0019_ sg13g2_dfrbpq_1
XFILLER_21_299 VPWR VGND sg13g2_decap_8
X_4668_ net671 net722 _0221_ VPWR VGND sg13g2_nor2_1
X_3619_ _1348_ VPWR _1349_ VGND _1312_ _1324_ sg13g2_o21ai_1
X_4770__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_1_616 VPWR VGND sg13g2_decap_8
X_4599_ net653 net704 _0152_ VPWR VGND sg13g2_nor2_1
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_48_108 VPWR VGND sg13g2_decap_8
XFILLER_29_311 VPWR VGND sg13g2_decap_4
XFILLER_45_804 VPWR VGND sg13g2_decap_4
XFILLER_29_344 VPWR VGND sg13g2_fill_1
XFILLER_29_355 VPWR VGND sg13g2_fill_1
XFILLER_17_528 VPWR VGND sg13g2_decap_8
XFILLER_44_347 VPWR VGND sg13g2_fill_2
XFILLER_44_358 VPWR VGND sg13g2_decap_8
XFILLER_13_701 VPWR VGND sg13g2_fill_2
XFILLER_12_211 VPWR VGND sg13g2_fill_2
XFILLER_40_531 VPWR VGND sg13g2_decap_8
XFILLER_8_215 VPWR VGND sg13g2_fill_1
XFILLER_12_299 VPWR VGND sg13g2_decap_8
XFILLER_5_911 VPWR VGND sg13g2_decap_8
XFILLER_5_26 VPWR VGND sg13g2_fill_2
XFILLER_5_988 VPWR VGND sg13g2_decap_8
XFILLER_47_185 VPWR VGND sg13g2_decap_4
X_3970_ _1682_ VPWR _1696_ VGND _1671_ _1677_ sg13g2_o21ai_1
X_4905__186 VPWR VGND net186 sg13g2_tiehi
X_2921_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\] net785 _0788_ _0283_
+ VPWR VGND sg13g2_mux2_1
X_2852_ _0775_ _0715_ _0773_ VPWR VGND sg13g2_nand2_2
X_2783_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[3\] net756 _0757_ _0464_
+ VPWR VGND sg13g2_mux2_1
X_4522_ net657 net708 _0075_ VPWR VGND sg13g2_nor2_1
X_4453_ net682 net733 _0008_ VPWR VGND sg13g2_nor2_1
X_3404_ _1134_ _1067_ _1132_ VPWR VGND sg13g2_xnor2_1
X_4384_ VGND VPWR _1993_ _2074_ _0624_ _2075_ sg13g2_a21oi_1
Xfanout706 net707 net706 VPWR VGND sg13g2_buf_8
Xfanout717 net718 net717 VPWR VGND sg13g2_buf_8
X_3335_ _1065_ _1060_ _1063_ VPWR VGND sg13g2_nand2_1
Xfanout728 net734 net728 VPWR VGND sg13g2_buf_8
Xfanout739 net745 net739 VPWR VGND sg13g2_buf_2
XFILLER_39_620 VPWR VGND sg13g2_decap_4
X_3266_ net749 _0997_ _0998_ _0368_ VPWR VGND sg13g2_nor3_1
X_5005_ net175 VGND VPWR _0552_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\]
+ _0200_ sg13g2_dfrbpq_1
XFILLER_38_163 VPWR VGND sg13g2_decap_8
X_3197_ _0951_ _0953_ _0954_ _0335_ VPWR VGND sg13g2_nor3_1
XFILLER_27_826 VPWR VGND sg13g2_fill_2
XFILLER_10_726 VPWR VGND sg13g2_decap_8
XFILLER_2_958 VPWR VGND sg13g2_decap_8
XFILLER_1_446 VPWR VGND sg13g2_decap_8
XFILLER_39_65 VPWR VGND sg13g2_fill_1
XFILLER_39_98 VPWR VGND sg13g2_decap_4
XFILLER_17_303 VPWR VGND sg13g2_fill_1
XFILLER_44_111 VPWR VGND sg13g2_decap_8
XFILLER_44_166 VPWR VGND sg13g2_decap_8
XFILLER_26_870 VPWR VGND sg13g2_fill_1
XFILLER_13_520 VPWR VGND sg13g2_decap_4
XFILLER_41_884 VPWR VGND sg13g2_fill_2
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_4_273 VPWR VGND sg13g2_fill_1
XFILLER_45_1024 VPWR VGND sg13g2_fill_1
XFILLER_45_1013 VPWR VGND sg13g2_decap_8
X_3120_ _0902_ _0797_ videogen.fancy_shader.video_x\[4\] VPWR VGND sg13g2_nand2b_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_49_995 VPWR VGND sg13g2_decap_8
X_3051_ net601 net602 _0842_ VPWR VGND sg13g2_xor2_1
XFILLER_24_807 VPWR VGND sg13g2_fill_1
X_4807__360 VPWR VGND net360 sg13g2_tiehi
XFILLER_35_166 VPWR VGND sg13g2_decap_8
X_3953_ _1678_ VPWR _1679_ VGND _1652_ _1656_ sg13g2_o21ai_1
X_2904_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\] _0785_ _0297_
+ VPWR VGND sg13g2_mux2_1
X_3884_ _1611_ _1612_ net612 _1613_ VPWR VGND sg13g2_nand3_1
X_2835_ _0728_ _0762_ _0770_ VPWR VGND sg13g2_nor2_2
X_2766_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\] _0753_ _0477_
+ VPWR VGND sg13g2_mux2_1
X_2697_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\] _0739_ _0541_
+ VPWR VGND sg13g2_mux2_1
X_4505_ net663 net724 _0058_ VPWR VGND sg13g2_nor2_1
X_4436_ _2126_ _1989_ _2125_ VPWR VGND sg13g2_nand2_1
X_4367_ VGND VPWR _2060_ _2061_ _0621_ net570 sg13g2_a21oi_1
X_3318_ _1028_ _1008_ _1048_ VPWR VGND sg13g2_nor2b_1
Xfanout547 _1176_ net547 VPWR VGND sg13g2_buf_8
Xfanout569 net571 net569 VPWR VGND sg13g2_buf_8
X_4298_ _2000_ net797 _1999_ VPWR VGND sg13g2_nand2b_1
Xfanout558 _1255_ net558 VPWR VGND sg13g2_buf_8
X_3249_ net748 _0987_ _0988_ _0361_ VPWR VGND sg13g2_nor3_1
X_5025__365 VPWR VGND net365 sg13g2_tiehi
XFILLER_39_472 VPWR VGND sg13g2_fill_2
XFILLER_26_111 VPWR VGND sg13g2_fill_2
XFILLER_42_604 VPWR VGND sg13g2_fill_1
XFILLER_26_133 VPWR VGND sg13g2_fill_1
XFILLER_23_840 VPWR VGND sg13g2_fill_2
XFILLER_41_55 VPWR VGND sg13g2_fill_1
XFILLER_41_44 VPWR VGND sg13g2_decap_8
X_4889__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_2_744 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_fill_1
XFILLER_49_247 VPWR VGND sg13g2_fill_1
XFILLER_2_49 VPWR VGND sg13g2_decap_8
X_4789__396 VPWR VGND net396 sg13g2_tiehi
XFILLER_46_921 VPWR VGND sg13g2_decap_8
XFILLER_18_623 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_fill_1
XFILLER_18_656 VPWR VGND sg13g2_decap_8
XFILLER_46_998 VPWR VGND sg13g2_decap_8
XFILLER_17_166 VPWR VGND sg13g2_decap_8
X_2620_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\] _0716_ _0595_
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_1023 VPWR VGND sg13g2_decap_4
X_2551_ videogen.fancy_shader.video_x\[8\] videogen.fancy_shader.video_x\[9\] _0666_
+ VPWR VGND sg13g2_nor2b_1
X_4221_ _1929_ tmds_red.n114 _1928_ VPWR VGND sg13g2_xnor2_1
X_4152_ _1874_ _1174_ _1875_ VPWR VGND sg13g2_xor2_1
X_4083_ _1806_ _1751_ _1805_ VPWR VGND sg13g2_xnor2_1
X_3103_ VGND VPWR tmds_red.n100 _0891_ _0274_ _0892_ sg13g2_a21oi_1
XFILLER_49_781 VPWR VGND sg13g2_fill_1
XFILLER_37_921 VPWR VGND sg13g2_decap_4
X_3034_ red_tmds_par\[9\] net696 serialize.n427\[9\] VPWR VGND sg13g2_and2_1
X_4985_ net258 VGND VPWR _0532_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\]
+ _0180_ sg13g2_dfrbpq_1
X_3936_ _1662_ _1657_ _1661_ VPWR VGND sg13g2_nand2_1
XFILLER_20_876 VPWR VGND sg13g2_decap_8
X_3867_ net597 _1595_ _1596_ VPWR VGND sg13g2_nor2_1
X_2818_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\] net778 _0766_ _0438_
+ VPWR VGND sg13g2_mux2_1
X_3798_ net616 VPWR _1528_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[3\]
+ net578 sg13g2_o21ai_1
X_2749_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\] net772 _0749_ _0490_
+ VPWR VGND sg13g2_mux2_1
X_4419_ _2109_ tmds_blue.dc_balancing_reg\[3\] _2080_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_921 VPWR VGND sg13g2_decap_8
XFILLER_43_935 VPWR VGND sg13g2_decap_8
XFILLER_42_401 VPWR VGND sg13g2_decap_8
XFILLER_27_464 VPWR VGND sg13g2_fill_2
XFILLER_27_486 VPWR VGND sg13g2_fill_1
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_42_456 VPWR VGND sg13g2_fill_2
XFILLER_35_1012 VPWR VGND sg13g2_decap_8
XFILLER_11_821 VPWR VGND sg13g2_fill_1
XFILLER_6_313 VPWR VGND sg13g2_decap_4
XFILLER_37_228 VPWR VGND sg13g2_decap_4
XFILLER_19_921 VPWR VGND sg13g2_decap_8
XFILLER_46_751 VPWR VGND sg13g2_fill_1
XFILLER_19_998 VPWR VGND sg13g2_decap_8
XFILLER_33_434 VPWR VGND sg13g2_fill_1
XFILLER_33_445 VPWR VGND sg13g2_fill_2
XFILLER_34_979 VPWR VGND sg13g2_decap_8
X_4770_ net62 VGND VPWR _0321_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\]
+ net631 sg13g2_dfrbpq_2
X_3721_ net749 net1 _1451_ VPWR VGND sg13g2_nor2_1
X_3652_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\] net559 _1382_ VPWR
+ VGND sg13g2_nor2_1
X_2603_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\] _0708_ _0604_
+ VPWR VGND sg13g2_mux2_1
X_3583_ net593 VPWR _1313_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\]
+ net562 sg13g2_o21ai_1
X_2534_ VPWR _0652_ tmds_red.dc_balancing_reg\[4\] VGND sg13g2_inv_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_4204_ VGND VPWR _0885_ _1916_ _1920_ _0647_ sg13g2_a21oi_1
X_4135_ _1798_ _1857_ _1858_ VPWR VGND sg13g2_nor2_1
XFILLER_28_217 VPWR VGND sg13g2_decap_8
X_4066_ _1789_ _1769_ _1788_ VPWR VGND sg13g2_xnor2_1
X_3017_ net440 green_tmds_par\[2\] net697 serialize.n428\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_25_913 VPWR VGND sg13g2_decap_8
X_4968_ net347 VGND VPWR _0515_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\]
+ _0163_ sg13g2_dfrbpq_1
X_3919_ _1637_ _1644_ _1645_ VPWR VGND sg13g2_and2_1
X_4899_ net198 VGND VPWR _0450_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\]
+ _0107_ sg13g2_dfrbpq_1
X_5059__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_3_327 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_fill_1
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_28_773 VPWR VGND sg13g2_fill_1
XFILLER_16_957 VPWR VGND sg13g2_decap_8
XFILLER_27_294 VPWR VGND sg13g2_fill_2
XFILLER_15_456 VPWR VGND sg13g2_fill_2
XFILLER_31_927 VPWR VGND sg13g2_decap_8
XFILLER_8_15 VPWR VGND sg13g2_fill_1
XFILLER_15_489 VPWR VGND sg13g2_fill_1
XFILLER_11_640 VPWR VGND sg13g2_decap_8
XFILLER_10_161 VPWR VGND sg13g2_decap_4
XFILLER_11_662 VPWR VGND sg13g2_decap_4
XFILLER_10_194 VPWR VGND sg13g2_decap_4
XFILLER_12_90 VPWR VGND sg13g2_decap_4
XFILLER_6_187 VPWR VGND sg13g2_decap_4
XFILLER_3_883 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_fill_2
XFILLER_34_710 VPWR VGND sg13g2_decap_8
XFILLER_18_294 VPWR VGND sg13g2_decap_8
XFILLER_19_795 VPWR VGND sg13g2_fill_2
XFILLER_22_949 VPWR VGND sg13g2_decap_8
X_4822_ net337 VGND VPWR _0373_ tmds_blue.n100 net640 sg13g2_dfrbpq_1
X_4753_ net86 VGND VPWR _0304_ videogen.fancy_shader.video_x\[1\] net636 sg13g2_dfrbpq_2
X_3704_ net594 _1428_ _1433_ _1434_ VPWR VGND sg13g2_nor3_1
XFILLER_30_993 VPWR VGND sg13g2_decap_8
X_4684_ net666 net717 _0237_ VPWR VGND sg13g2_nor2_1
X_3635_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\] net585 _1365_ VPWR
+ VGND sg13g2_nor2_1
X_4915__166 VPWR VGND net166 sg13g2_tiehi
X_3566_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\] net580 _1296_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_3497_ _1227_ net545 _1225_ VPWR VGND sg13g2_xnor2_1
X_2517_ VPWR _0635_ videogen.fancy_shader.n646\[0\] VGND sg13g2_inv_1
X_4731__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_25_1011 VPWR VGND sg13g2_decap_8
X_5098_ net801 VGND VPWR serialize.n431\[3\] serialize.n420\[1\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4118_ _1797_ _1031_ _1841_ VPWR VGND sg13g2_xor2_1
XFILLER_37_570 VPWR VGND sg13g2_fill_1
X_4049_ _1626_ net546 _1772_ VPWR VGND sg13g2_xor2_1
XFILLER_13_916 VPWR VGND sg13g2_decap_8
XFILLER_40_779 VPWR VGND sg13g2_fill_1
XFILLER_8_408 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_fill_2
XFILLER_32_1004 VPWR VGND sg13g2_decap_8
XFILLER_21_971 VPWR VGND sg13g2_decap_8
XFILLER_20_481 VPWR VGND sg13g2_fill_2
XFILLER_0_842 VPWR VGND sg13g2_decap_8
Xhold8 serialize.bit_cnt\[0\] VPWR VGND net413 sg13g2_dlygate4sd3_1
XFILLER_47_334 VPWR VGND sg13g2_decap_8
XFILLER_47_389 VPWR VGND sg13g2_fill_1
X_5040__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_16_721 VPWR VGND sg13g2_decap_8
XFILLER_16_765 VPWR VGND sg13g2_decap_4
XFILLER_15_275 VPWR VGND sg13g2_decap_8
XFILLER_15_286 VPWR VGND sg13g2_fill_2
XFILLER_30_212 VPWR VGND sg13g2_fill_1
XFILLER_12_960 VPWR VGND sg13g2_decap_8
XFILLER_30_256 VPWR VGND sg13g2_fill_1
XFILLER_8_975 VPWR VGND sg13g2_decap_8
XFILLER_7_474 VPWR VGND sg13g2_fill_2
XFILLER_48_1000 VPWR VGND sg13g2_decap_8
X_3420_ _1127_ _1133_ _1149_ _1150_ VPWR VGND sg13g2_or3_1
X_4951__399 VPWR VGND net399 sg13g2_tiehi
X_3351_ videogen.fancy_shader.video_y\[6\] videogen.fancy_shader.n646\[6\] _1081_
+ VPWR VGND sg13g2_and2_1
X_3282_ _1012_ videogen.fancy_shader.n646\[0\] net630 VPWR VGND sg13g2_nand2_1
X_5021_ net43 VGND VPWR _0568_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\]
+ _0216_ sg13g2_dfrbpq_1
XFILLER_39_879 VPWR VGND sg13g2_fill_1
XFILLER_39_868 VPWR VGND sg13g2_fill_2
XFILLER_26_529 VPWR VGND sg13g2_decap_8
XFILLER_0_71 VPWR VGND sg13g2_fill_1
XFILLER_0_60 VPWR VGND sg13g2_decap_8
XFILLER_0_1024 VPWR VGND sg13g2_decap_4
XFILLER_19_581 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_fill_2
XFILLER_21_212 VPWR VGND sg13g2_decap_8
XFILLER_10_919 VPWR VGND sg13g2_decap_8
X_4805_ net364 VGND VPWR _0356_ videogen.fancy_shader.video_y\[0\] net637 sg13g2_dfrbpq_2
XFILLER_22_768 VPWR VGND sg13g2_decap_8
X_2997_ net699 net409 serialize.n431\[0\] VPWR VGND sg13g2_nor2b_1
XFILLER_9_91 VPWR VGND sg13g2_fill_2
X_4736_ net119 VGND VPWR _0287_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\]
+ _0018_ sg13g2_dfrbpq_1
X_4667_ net686 net737 _0220_ VPWR VGND sg13g2_nor2_1
X_3618_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1347_ _1348_ VPWR VGND
+ sg13g2_nor2_1
X_4598_ net653 net704 _0151_ VPWR VGND sg13g2_nor2_1
XFILLER_0_116 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_fill_1
X_3549_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\] net553 _1279_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_149 VPWR VGND sg13g2_decap_8
X_4967__351 VPWR VGND net351 sg13g2_tiehi
X_5078__31 VPWR VGND net31 sg13g2_tiehi
XFILLER_44_326 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_fill_2
XFILLER_29_389 VPWR VGND sg13g2_decap_8
XFILLER_13_713 VPWR VGND sg13g2_decap_8
X_4974__300 VPWR VGND net300 sg13g2_tiehi
XFILLER_12_245 VPWR VGND sg13g2_decap_8
XFILLER_8_227 VPWR VGND sg13g2_decap_4
XFILLER_8_205 VPWR VGND sg13g2_decap_4
XFILLER_5_967 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_5_38 VPWR VGND sg13g2_decap_8
XFILLER_29_890 VPWR VGND sg13g2_decap_8
X_2920_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\] net776 _0788_ _0284_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_510 VPWR VGND sg13g2_fill_2
X_2851_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\] _0774_ _0413_
+ VPWR VGND sg13g2_mux2_1
X_4799__376 VPWR VGND net376 sg13g2_tiehi
X_2782_ _0723_ _0751_ _0757_ VPWR VGND sg13g2_nor2b_2
X_4521_ net658 net709 _0074_ VPWR VGND sg13g2_nor2_1
X_4452_ net680 net731 _0007_ VPWR VGND sg13g2_nor2_1
X_3403_ _1067_ _1132_ _1133_ VPWR VGND sg13g2_nor2_1
X_4383_ _0836_ VPWR _2075_ VGND _1993_ _2074_ sg13g2_o21ai_1
Xfanout718 net724 net718 VPWR VGND sg13g2_buf_8
X_3334_ VGND VPWR _1064_ _1063_ _1060_ sg13g2_or2_1
Xfanout707 net746 net707 VPWR VGND sg13g2_buf_8
Xfanout729 net734 net729 VPWR VGND sg13g2_buf_1
X_3265_ _0998_ videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ videogen.test_lut_thingy.gol_counter_reg\[2\] VPWR VGND sg13g2_and3_1
X_5004_ net179 VGND VPWR _0551_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\]
+ _0199_ sg13g2_dfrbpq_1
X_3196_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\] _0802_ _0954_ VPWR
+ VGND sg13g2_and2_1
XFILLER_22_576 VPWR VGND sg13g2_decap_8
XFILLER_10_749 VPWR VGND sg13g2_decap_8
X_4719_ net145 VGND VPWR _0270_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\]
+ _0009_ sg13g2_dfrbpq_1
XFILLER_30_79 VPWR VGND sg13g2_fill_1
XFILLER_2_937 VPWR VGND sg13g2_decap_8
XFILLER_1_414 VPWR VGND sg13g2_fill_1
XFILLER_39_88 VPWR VGND sg13g2_fill_1
XFILLER_18_827 VPWR VGND sg13g2_fill_1
XFILLER_29_175 VPWR VGND sg13g2_fill_2
XFILLER_38_1021 VPWR VGND sg13g2_decap_8
XFILLER_32_329 VPWR VGND sg13g2_fill_2
XFILLER_9_536 VPWR VGND sg13g2_fill_2
XFILLER_9_569 VPWR VGND sg13g2_fill_1
XFILLER_5_742 VPWR VGND sg13g2_decap_4
XFILLER_4_285 VPWR VGND sg13g2_decap_8
XFILLER_20_90 VPWR VGND sg13g2_decap_8
X_3050_ _0841_ net602 net601 VPWR VGND sg13g2_nand2b_1
XFILLER_49_974 VPWR VGND sg13g2_decap_8
XFILLER_36_657 VPWR VGND sg13g2_fill_2
XFILLER_17_860 VPWR VGND sg13g2_fill_1
X_3952_ _1651_ VPWR _1678_ VGND _1635_ _1656_ sg13g2_o21ai_1
X_2903_ net753 videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\] _0785_ _0298_
+ VPWR VGND sg13g2_mux2_1
X_3883_ net598 VPWR _1612_ VGND _1556_ _1561_ sg13g2_o21ai_1
X_2834_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\] net783 _0769_ _0425_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_395 VPWR VGND sg13g2_decap_4
X_4504_ net651 net702 _0057_ VPWR VGND sg13g2_nor2_1
X_2765_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\] _0753_ _0478_
+ VPWR VGND sg13g2_mux2_1
X_2696_ _0739_ _0698_ _0731_ VPWR VGND sg13g2_nand2_2
X_4435_ _2125_ _2123_ _2124_ _2122_ _1991_ VPWR VGND sg13g2_a22oi_1
X_4366_ VGND VPWR _0847_ _2055_ _2061_ _0840_ sg13g2_a21oi_1
X_3317_ _1009_ _1029_ _1047_ VPWR VGND sg13g2_and2_1
Xfanout548 _0855_ net548 VPWR VGND sg13g2_buf_8
X_4297_ net606 hsync _1999_ VPWR VGND sg13g2_nor2b_1
Xfanout559 net568 net559 VPWR VGND sg13g2_buf_8
X_3248_ _0988_ videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.video_y\[4\]
+ _0984_ VPWR VGND sg13g2_and3_2
X_3179_ _0943_ _0636_ _0941_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_624 VPWR VGND sg13g2_fill_1
XFILLER_15_819 VPWR VGND sg13g2_decap_4
XFILLER_27_679 VPWR VGND sg13g2_fill_1
XFILLER_42_627 VPWR VGND sg13g2_decap_4
XFILLER_42_649 VPWR VGND sg13g2_fill_1
XFILLER_41_148 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_fill_1
XFILLER_41_159 VPWR VGND sg13g2_fill_1
XFILLER_23_885 VPWR VGND sg13g2_decap_8
XFILLER_22_384 VPWR VGND sg13g2_decap_4
XFILLER_2_723 VPWR VGND sg13g2_decap_4
XFILLER_29_1009 VPWR VGND sg13g2_decap_8
XFILLER_1_288 VPWR VGND sg13g2_fill_2
XFILLER_49_259 VPWR VGND sg13g2_fill_2
XFILLER_46_900 VPWR VGND sg13g2_decap_8
XFILLER_46_977 VPWR VGND sg13g2_decap_8
XFILLER_17_123 VPWR VGND sg13g2_decap_8
XFILLER_17_134 VPWR VGND sg13g2_fill_2
XFILLER_32_148 VPWR VGND sg13g2_fill_1
XFILLER_9_311 VPWR VGND sg13g2_fill_1
XFILLER_13_384 VPWR VGND sg13g2_decap_8
XFILLER_12_1002 VPWR VGND sg13g2_decap_8
X_2550_ _0662_ _0664_ _0665_ VPWR VGND sg13g2_nor2b_2
X_4220_ _1928_ tmds_red.n132 tmds_red.dc_balancing_reg\[1\] VPWR VGND sg13g2_xnor2_1
X_4151_ _1874_ _1725_ _1873_ VPWR VGND sg13g2_nand2_1
X_4082_ _1801_ _1063_ _1805_ VPWR VGND sg13g2_xor2_1
X_3102_ _0836_ VPWR _0892_ VGND tmds_red.n100 _0891_ sg13g2_o21ai_1
X_3033_ red_tmds_par\[8\] net696 serialize.n427\[8\] VPWR VGND sg13g2_and2_1
XFILLER_23_126 VPWR VGND sg13g2_decap_8
X_4984_ net262 VGND VPWR _0531_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\]
+ _0179_ sg13g2_dfrbpq_1
X_3935_ _1651_ _1659_ _1661_ VPWR VGND sg13g2_nor2_1
X_3866_ net621 _1594_ _1595_ VPWR VGND sg13g2_nor2_1
XFILLER_20_844 VPWR VGND sg13g2_fill_2
X_3797_ _1523_ _1524_ _1525_ _1526_ _1527_ VPWR VGND sg13g2_nor4_1
X_2817_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\] net767 _0766_ _0439_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_899 VPWR VGND sg13g2_fill_1
X_2748_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\] net762 _0749_ _0491_
+ VPWR VGND sg13g2_mux2_1
X_4418_ _2081_ VPWR _2108_ VGND _2080_ _2107_ sg13g2_o21ai_1
X_2679_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\] _0735_ _0555_
+ VPWR VGND sg13g2_mux2_1
X_4349_ _2044_ _2026_ _2028_ VPWR VGND sg13g2_nand2_1
XFILLER_28_900 VPWR VGND sg13g2_decap_8
XFILLER_27_410 VPWR VGND sg13g2_fill_2
X_4925__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_42_435 VPWR VGND sg13g2_fill_2
X_4741__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_10_343 VPWR VGND sg13g2_fill_2
XFILLER_7_859 VPWR VGND sg13g2_fill_2
XFILLER_7_826 VPWR VGND sg13g2_decap_4
X_5071__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_7_0 VPWR VGND sg13g2_decap_4
XFILLER_2_564 VPWR VGND sg13g2_decap_4
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_977 VPWR VGND sg13g2_decap_8
XFILLER_46_796 VPWR VGND sg13g2_decap_8
XFILLER_18_476 VPWR VGND sg13g2_decap_4
XFILLER_20_129 VPWR VGND sg13g2_decap_8
X_3720_ _1450_ _1352_ _1449_ VPWR VGND sg13g2_nand2_1
XFILLER_9_141 VPWR VGND sg13g2_fill_2
XFILLER_9_174 VPWR VGND sg13g2_decap_8
X_3651_ net596 VPWR _1381_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\]
+ net583 sg13g2_o21ai_1
X_2602_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\] _0708_ _0605_
+ VPWR VGND sg13g2_mux2_1
X_3582_ net618 _1306_ _1311_ _1312_ VPWR VGND sg13g2_nor3_1
X_2533_ VPWR _0651_ videogen.test_lut_thingy.gol_counter_reg\[2\] VGND sg13g2_inv_1
X_4203_ VPWR _1919_ _1918_ VGND sg13g2_inv_1
XFILLER_3_60 VPWR VGND sg13g2_fill_2
X_4134_ _1857_ _1854_ _1855_ VPWR VGND sg13g2_nand2_1
X_4065_ VGND VPWR _1773_ _1776_ _1788_ _1787_ sg13g2_a21oi_1
X_3016_ _0834_ VPWR serialize.n428\[1\] VGND _0655_ net700 sg13g2_o21ai_1
XFILLER_36_251 VPWR VGND sg13g2_fill_1
XFILLER_25_969 VPWR VGND sg13g2_decap_8
XFILLER_12_608 VPWR VGND sg13g2_decap_4
XFILLER_19_1019 VPWR VGND sg13g2_decap_4
XFILLER_24_457 VPWR VGND sg13g2_fill_1
X_4967_ net351 VGND VPWR _0514_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\]
+ _0162_ sg13g2_dfrbpq_1
X_3918_ _1640_ _1641_ _1643_ _1644_ VPWR VGND sg13g2_or3_1
X_4898_ net200 VGND VPWR _0449_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\]
+ _0106_ sg13g2_dfrbpq_1
X_3849_ net595 VPWR _1578_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\]
+ net567 sg13g2_o21ai_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_218 VPWR VGND sg13g2_decap_8
XFILLER_28_741 VPWR VGND sg13g2_decap_8
XFILLER_27_240 VPWR VGND sg13g2_fill_2
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_15_435 VPWR VGND sg13g2_decap_8
XFILLER_16_936 VPWR VGND sg13g2_decap_8
XFILLER_31_906 VPWR VGND sg13g2_decap_8
XFILLER_7_612 VPWR VGND sg13g2_fill_1
XFILLER_3_862 VPWR VGND sg13g2_decap_8
XFILLER_18_251 VPWR VGND sg13g2_decap_8
XFILLER_19_763 VPWR VGND sg13g2_decap_4
XFILLER_18_262 VPWR VGND sg13g2_fill_2
XFILLER_33_254 VPWR VGND sg13g2_decap_4
X_4821_ net338 VGND VPWR _0372_ tmds_blue.n193 net641 sg13g2_dfrbpq_2
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_22_928 VPWR VGND sg13g2_decap_8
X_4752_ net87 VGND VPWR _0303_ videogen.fancy_shader.video_x\[0\] net638 sg13g2_dfrbpq_2
XFILLER_21_449 VPWR VGND sg13g2_decap_8
X_3703_ _1429_ _1430_ _1431_ _1432_ _1433_ VPWR VGND sg13g2_nor4_1
XFILLER_30_972 VPWR VGND sg13g2_decap_8
X_4683_ net668 net714 _0236_ VPWR VGND sg13g2_nor2_1
X_3634_ net615 VPWR _1364_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\]
+ net562 sg13g2_o21ai_1
X_3565_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\] net556 _1295_ VPWR
+ VGND sg13g2_nor2_1
X_2516_ VPWR _0634_ videogen.fancy_shader.n646\[5\] VGND sg13g2_inv_1
X_3496_ _1226_ net545 _1225_ VPWR VGND sg13g2_nand2_1
X_5097_ net801 VGND VPWR serialize.n431\[2\] serialize.n420\[0\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4117_ _1840_ _1802_ _1837_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_538 VPWR VGND sg13g2_decap_8
X_4048_ _1727_ VPWR _1771_ VGND _1027_ _1770_ sg13g2_o21ai_1
XFILLER_17_25 VPWR VGND sg13g2_fill_1
XFILLER_37_593 VPWR VGND sg13g2_decap_4
XFILLER_33_13 VPWR VGND sg13g2_fill_1
XFILLER_21_950 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_0_821 VPWR VGND sg13g2_decap_8
Xhold9 serialize.n414\[3\] VPWR VGND net414 sg13g2_dlygate4sd3_1
XFILLER_0_898 VPWR VGND sg13g2_decap_8
XFILLER_47_379 VPWR VGND sg13g2_decap_4
XFILLER_28_560 VPWR VGND sg13g2_fill_2
XFILLER_35_519 VPWR VGND sg13g2_fill_2
XFILLER_43_541 VPWR VGND sg13g2_decap_4
XFILLER_15_243 VPWR VGND sg13g2_fill_2
XFILLER_16_744 VPWR VGND sg13g2_decap_8
XFILLER_30_202 VPWR VGND sg13g2_fill_2
XFILLER_31_747 VPWR VGND sg13g2_decap_8
XFILLER_8_954 VPWR VGND sg13g2_decap_8
XFILLER_7_442 VPWR VGND sg13g2_fill_1
XFILLER_11_493 VPWR VGND sg13g2_decap_4
XFILLER_23_90 VPWR VGND sg13g2_fill_1
X_3350_ _1079_ VPWR _1080_ VGND _1049_ _1077_ sg13g2_o21ai_1
XFILLER_3_670 VPWR VGND sg13g2_decap_8
X_3281_ _1011_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_x\[1\]
+ VPWR VGND sg13g2_nand2_1
X_5020_ net51 VGND VPWR _0567_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\]
+ _0215_ sg13g2_dfrbpq_1
XFILLER_38_313 VPWR VGND sg13g2_decap_8
XFILLER_0_1003 VPWR VGND sg13g2_decap_8
XFILLER_34_585 VPWR VGND sg13g2_fill_2
X_4804_ net366 VGND VPWR _0355_ videogen.fancy_shader.n646\[9\] net633 sg13g2_dfrbpq_2
X_2996_ net413 net695 serialize.n433\[0\] VPWR VGND sg13g2_nor2_1
X_4735_ net121 VGND VPWR _0286_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\]
+ _0017_ sg13g2_dfrbpq_1
X_4666_ net671 net722 _0219_ VPWR VGND sg13g2_nor2_1
X_4597_ net654 net705 _0150_ VPWR VGND sg13g2_nor2_1
X_3617_ net612 _1335_ _1346_ _1347_ VPWR VGND sg13g2_nor3_1
X_3548_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\] net563 _1278_ VPWR
+ VGND sg13g2_nor2_1
X_3479_ _1197_ VPWR _1209_ VGND _1205_ _1208_ sg13g2_o21ai_1
XFILLER_29_335 VPWR VGND sg13g2_decap_8
XFILLER_28_68 VPWR VGND sg13g2_decap_4
XFILLER_44_349 VPWR VGND sg13g2_fill_1
XFILLER_40_500 VPWR VGND sg13g2_decap_4
XFILLER_12_213 VPWR VGND sg13g2_fill_1
XFILLER_12_224 VPWR VGND sg13g2_fill_2
XFILLER_13_769 VPWR VGND sg13g2_fill_2
XFILLER_40_566 VPWR VGND sg13g2_decap_8
XFILLER_12_257 VPWR VGND sg13g2_fill_2
XFILLER_40_599 VPWR VGND sg13g2_fill_1
XFILLER_5_946 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_4
XFILLER_48_611 VPWR VGND sg13g2_decap_8
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_48_655 VPWR VGND sg13g2_decap_8
XFILLER_44_883 VPWR VGND sg13g2_decap_8
X_2850_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\] _0774_ _0414_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
X_2781_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\] _0756_ _0465_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_762 VPWR VGND sg13g2_fill_2
XFILLER_8_751 VPWR VGND sg13g2_decap_8
X_4520_ net678 net726 _0073_ VPWR VGND sg13g2_nor2_1
X_4451_ VGND VPWR _2121_ _2139_ _0627_ net571 sg13g2_a21oi_1
XFILLER_8_795 VPWR VGND sg13g2_decap_4
X_3402_ VGND VPWR _1128_ _1130_ _1132_ _1131_ sg13g2_a21oi_1
X_4382_ _2074_ tmds_blue.n132 _2073_ VPWR VGND sg13g2_xnor2_1
X_3333_ _1063_ _1061_ _1062_ VPWR VGND sg13g2_xnor2_1
Xfanout708 net711 net708 VPWR VGND sg13g2_buf_8
Xfanout719 net720 net719 VPWR VGND sg13g2_buf_8
XFILLER_39_600 VPWR VGND sg13g2_fill_2
X_3264_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ _0997_ videogen.test_lut_thingy.gol_counter_reg\[2\] sg13g2_a21oi_1
X_5003_ net183 VGND VPWR _0550_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\]
+ _0198_ sg13g2_dfrbpq_1
XFILLER_39_666 VPWR VGND sg13g2_decap_8
X_3195_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\] _0802_ _0953_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_22_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_806 VPWR VGND sg13g2_decap_8
XFILLER_27_828 VPWR VGND sg13g2_fill_1
XFILLER_39_699 VPWR VGND sg13g2_fill_1
XFILLER_26_316 VPWR VGND sg13g2_fill_2
XFILLER_35_883 VPWR VGND sg13g2_fill_2
XFILLER_14_37 VPWR VGND sg13g2_fill_2
XFILLER_14_59 VPWR VGND sg13g2_decap_8
XFILLER_22_555 VPWR VGND sg13g2_decap_8
X_2979_ _0825_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\]
+ _0822_ VPWR VGND sg13g2_and3_2
X_4718_ net147 VGND VPWR _0269_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\]
+ _0008_ sg13g2_dfrbpq_1
X_4649_ net659 net710 _0202_ VPWR VGND sg13g2_nor2_1
XFILLER_2_916 VPWR VGND sg13g2_decap_8
XFILLER_39_23 VPWR VGND sg13g2_decap_8
XFILLER_49_419 VPWR VGND sg13g2_decap_8
XFILLER_49_408 VPWR VGND sg13g2_decap_8
XFILLER_39_34 VPWR VGND sg13g2_fill_2
XFILLER_45_625 VPWR VGND sg13g2_decap_8
XFILLER_18_839 VPWR VGND sg13g2_decap_8
XFILLER_38_1000 VPWR VGND sg13g2_decap_8
XFILLER_25_393 VPWR VGND sg13g2_decap_4
XFILLER_41_886 VPWR VGND sg13g2_fill_1
XFILLER_40_341 VPWR VGND sg13g2_fill_1
XFILLER_9_526 VPWR VGND sg13g2_fill_2
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_5_787 VPWR VGND sg13g2_decap_8
XFILLER_49_953 VPWR VGND sg13g2_decap_8
XFILLER_1_993 VPWR VGND sg13g2_decap_8
XFILLER_35_102 VPWR VGND sg13g2_fill_1
X_3951_ _1677_ _1672_ _1674_ _1676_ VPWR VGND sg13g2_and3_1
XFILLER_17_883 VPWR VGND sg13g2_decap_8
XFILLER_44_691 VPWR VGND sg13g2_decap_8
XFILLER_44_680 VPWR VGND sg13g2_fill_1
XFILLER_17_894 VPWR VGND sg13g2_fill_2
X_2902_ _0785_ _0720_ _0727_ VPWR VGND sg13g2_nand2_2
X_3882_ _1607_ _1610_ net615 _1611_ VPWR VGND sg13g2_nand3_1
X_2833_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\] net773 _0769_ _0426_
+ VPWR VGND sg13g2_mux2_1
X_2764_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\] _0753_ _0479_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_592 VPWR VGND sg13g2_fill_1
X_4503_ net652 net703 _0056_ VPWR VGND sg13g2_nor2_1
X_2695_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\] _0738_ _0542_
+ VPWR VGND sg13g2_mux2_1
X_4434_ VGND VPWR _2102_ _2113_ _2124_ _1991_ sg13g2_a21oi_1
X_4365_ _2060_ _2059_ _0847_ VPWR VGND sg13g2_nand2b_1
X_3316_ _1046_ _1041_ _1044_ VPWR VGND sg13g2_xnor2_1
X_4296_ _1994_ _1998_ _0611_ VPWR VGND sg13g2_nor2_1
Xfanout549 net558 net549 VPWR VGND sg13g2_buf_8
XFILLER_39_441 VPWR VGND sg13g2_fill_1
X_3247_ videogen.fancy_shader.video_y\[5\] _0985_ _0987_ VPWR VGND sg13g2_nor2_1
XFILLER_39_496 VPWR VGND sg13g2_decap_4
X_3178_ _0940_ _0942_ _0328_ VPWR VGND sg13g2_nor2_1
XFILLER_26_124 VPWR VGND sg13g2_decap_8
XFILLER_23_842 VPWR VGND sg13g2_fill_1
XFILLER_10_525 VPWR VGND sg13g2_fill_2
X_4936__402 VPWR VGND net402 sg13g2_tiehi
X_4858__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_2_702 VPWR VGND sg13g2_fill_1
XFILLER_9_4 VPWR VGND sg13g2_fill_2
XFILLER_1_267 VPWR VGND sg13g2_decap_8
XFILLER_17_102 VPWR VGND sg13g2_decap_8
XFILLER_46_956 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_9_301 VPWR VGND sg13g2_decap_4
XFILLER_14_853 VPWR VGND sg13g2_fill_1
XFILLER_41_672 VPWR VGND sg13g2_decap_8
XFILLER_14_886 VPWR VGND sg13g2_decap_8
XFILLER_15_91 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
X_4837__322 VPWR VGND net322 sg13g2_tiehi
X_4150_ _1873_ _1724_ _1175_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_790 VPWR VGND sg13g2_decap_8
X_3101_ VGND VPWR _0885_ _0891_ _0889_ _0884_ sg13g2_a21oi_2
X_4081_ _1063_ _1799_ _1052_ _1804_ VPWR VGND sg13g2_nand3_1
XFILLER_49_772 VPWR VGND sg13g2_decap_8
X_3032_ net424 red_tmds_par\[7\] net697 serialize.n427\[7\] VPWR VGND sg13g2_mux2_1
XFILLER_36_400 VPWR VGND sg13g2_fill_1
XFILLER_36_444 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_8
XFILLER_23_105 VPWR VGND sg13g2_decap_8
X_4983_ net266 VGND VPWR _0530_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\]
+ _0178_ sg13g2_dfrbpq_1
X_3934_ VPWR _1660_ _1659_ VGND sg13g2_inv_1
X_3865_ net625 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\] videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\]
+ net628 _1594_ VPWR VGND sg13g2_mux4_1
XFILLER_32_661 VPWR VGND sg13g2_decap_8
X_2816_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\] net757 _0766_ _0440_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_171 VPWR VGND sg13g2_decap_8
XFILLER_31_193 VPWR VGND sg13g2_fill_1
X_3796_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\] net556 _1526_ VPWR
+ VGND sg13g2_nor2_1
X_2747_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\] net752 _0749_ _0492_
+ VPWR VGND sg13g2_mux2_1
X_2678_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\] _0735_ _0556_
+ VPWR VGND sg13g2_mux2_1
X_4417_ VPWR _2107_ _2106_ VGND sg13g2_inv_1
X_4888__220 VPWR VGND net220 sg13g2_tiehi
X_4348_ VPWR _2043_ _2042_ VGND sg13g2_inv_1
XFILLER_47_709 VPWR VGND sg13g2_fill_2
X_4279_ VGND VPWR _1970_ _1982_ _1984_ _1983_ sg13g2_a21oi_1
XFILLER_39_260 VPWR VGND sg13g2_decap_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_23_672 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_fill_1
XFILLER_10_322 VPWR VGND sg13g2_fill_1
XFILLER_22_182 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_fill_2
XFILLER_10_377 VPWR VGND sg13g2_fill_2
XFILLER_2_532 VPWR VGND sg13g2_fill_2
XFILLER_42_1007 VPWR VGND sg13g2_decap_8
XFILLER_38_709 VPWR VGND sg13g2_fill_2
XFILLER_18_422 VPWR VGND sg13g2_fill_2
XFILLER_19_956 VPWR VGND sg13g2_decap_8
XFILLER_46_775 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_fill_2
XFILLER_20_108 VPWR VGND sg13g2_fill_1
XFILLER_13_171 VPWR VGND sg13g2_fill_1
X_3650_ _1376_ _1377_ _1378_ _1379_ _1380_ VPWR VGND sg13g2_nor4_1
X_2601_ _0708_ _0698_ _0706_ VPWR VGND sg13g2_nand2_2
X_3581_ _1307_ _1308_ _1309_ _1310_ _1311_ VPWR VGND sg13g2_nor4_1
X_2532_ VPWR _0650_ net2 VGND sg13g2_inv_1
XFILLER_6_893 VPWR VGND sg13g2_decap_8
XFILLER_5_370 VPWR VGND sg13g2_fill_1
X_4202_ VGND VPWR _1918_ _0884_ net548 sg13g2_or2_1
X_4133_ _1854_ _1855_ _1856_ VPWR VGND sg13g2_and2_1
X_4064_ VGND VPWR _1769_ _1782_ _1787_ _1780_ sg13g2_a21oi_1
X_5009__159 VPWR VGND net159 sg13g2_tiehi
X_3015_ _0834_ green_tmds_par\[1\] net698 VPWR VGND sg13g2_nand2_1
XFILLER_37_720 VPWR VGND sg13g2_fill_2
XFILLER_3_1023 VPWR VGND sg13g2_decap_4
XFILLER_36_230 VPWR VGND sg13g2_fill_1
XFILLER_24_425 VPWR VGND sg13g2_fill_1
XFILLER_25_948 VPWR VGND sg13g2_decap_8
XFILLER_36_285 VPWR VGND sg13g2_decap_8
X_4966_ net355 VGND VPWR _0513_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\]
+ _0161_ sg13g2_dfrbpq_1
XFILLER_11_108 VPWR VGND sg13g2_fill_1
X_4777__48 VPWR VGND net48 sg13g2_tiehi
X_4897_ net202 VGND VPWR _0448_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\]
+ _0105_ sg13g2_dfrbpq_1
X_3917_ _1642_ _1120_ _1643_ VPWR VGND sg13g2_xor2_1
X_3848_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\] net556 _1577_ VPWR
+ VGND sg13g2_nor2_1
X_3779_ _1505_ _1506_ _1507_ _1508_ _1509_ VPWR VGND sg13g2_nor4_1
XFILLER_22_59 VPWR VGND sg13g2_decap_8
XFILLER_3_307 VPWR VGND sg13g2_decap_4
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_27_252 VPWR VGND sg13g2_decap_8
X_4827__332 VPWR VGND net332 sg13g2_tiehi
XFILLER_15_458 VPWR VGND sg13g2_fill_1
XFILLER_24_981 VPWR VGND sg13g2_decap_8
XFILLER_30_417 VPWR VGND sg13g2_fill_2
XFILLER_8_39 VPWR VGND sg13g2_decap_4
XFILLER_11_631 VPWR VGND sg13g2_decap_4
XFILLER_30_439 VPWR VGND sg13g2_fill_2
X_4834__325 VPWR VGND net325 sg13g2_tiehi
XFILLER_40_9 VPWR VGND sg13g2_decap_4
XFILLER_3_852 VPWR VGND sg13g2_fill_1
XFILLER_3_841 VPWR VGND sg13g2_decap_8
XFILLER_46_594 VPWR VGND sg13g2_fill_1
XFILLER_33_211 VPWR VGND sg13g2_decap_4
XFILLER_22_907 VPWR VGND sg13g2_decap_8
X_4820_ net339 VGND VPWR _0371_ display_enable net640 sg13g2_dfrbpq_1
XFILLER_34_745 VPWR VGND sg13g2_decap_8
XFILLER_21_417 VPWR VGND sg13g2_decap_8
XFILLER_21_428 VPWR VGND sg13g2_fill_2
X_4751_ net89 VGND VPWR _0302_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\]
+ _0033_ sg13g2_dfrbpq_1
XFILLER_30_951 VPWR VGND sg13g2_decap_8
X_4682_ net664 net715 _0235_ VPWR VGND sg13g2_nor2_1
X_3702_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\] net586 _1432_ VPWR
+ VGND sg13g2_nor2_1
X_3633_ net622 _1357_ _1362_ _1363_ VPWR VGND sg13g2_nor3_1
X_3564_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\] net589 _1294_ VPWR
+ VGND sg13g2_nor2_1
X_2515_ VPWR _0633_ videogen.fancy_shader.video_y\[5\] VGND sg13g2_inv_1
X_3495_ _1223_ _1224_ _1225_ VPWR VGND _1221_ sg13g2_nand3b_1
X_4116_ _1839_ _1803_ _1837_ VPWR VGND sg13g2_xnor2_1
X_5096_ net801 VGND VPWR serialize.n431\[1\] serialize.n461 clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_44_509 VPWR VGND sg13g2_fill_2
X_4047_ _1018_ _1725_ _1770_ VPWR VGND sg13g2_nor2_1
XFILLER_24_233 VPWR VGND sg13g2_decap_8
XFILLER_24_244 VPWR VGND sg13g2_fill_2
XFILLER_12_406 VPWR VGND sg13g2_fill_2
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_12_439 VPWR VGND sg13g2_fill_2
X_4949_ net33 VGND VPWR _0496_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\]
+ _0153_ sg13g2_dfrbpq_1
X_4758__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_20_483 VPWR VGND sg13g2_fill_1
XFILLER_4_616 VPWR VGND sg13g2_decap_8
XFILLER_3_115 VPWR VGND sg13g2_fill_2
XFILLER_3_104 VPWR VGND sg13g2_fill_1
XFILLER_0_800 VPWR VGND sg13g2_decap_8
XFILLER_0_877 VPWR VGND sg13g2_decap_8
XFILLER_47_358 VPWR VGND sg13g2_decap_8
XFILLER_28_550 VPWR VGND sg13g2_fill_2
XFILLER_16_789 VPWR VGND sg13g2_decap_8
XFILLER_43_597 VPWR VGND sg13g2_decap_8
XFILLER_8_933 VPWR VGND sg13g2_decap_8
XFILLER_12_995 VPWR VGND sg13g2_decap_8
X_4764__73 VPWR VGND net73 sg13g2_tiehi
X_3280_ _1010_ _1007_ _1009_ VPWR VGND sg13g2_xnor2_1
X_4730__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_2_192 VPWR VGND sg13g2_decap_8
XFILLER_31_5 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_38_336 VPWR VGND sg13g2_fill_2
XFILLER_47_892 VPWR VGND sg13g2_decap_8
XFILLER_19_572 VPWR VGND sg13g2_decap_4
XFILLER_0_95 VPWR VGND sg13g2_decap_4
XFILLER_22_715 VPWR VGND sg13g2_decap_8
X_4803_ net368 VGND VPWR _0354_ videogen.fancy_shader.n646\[8\] net633 sg13g2_dfrbpq_1
X_4734_ net123 VGND VPWR _0285_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\]
+ _0016_ sg13g2_dfrbpq_1
X_2995_ serialize.n452 serialize.n450 clknet_1_1__leaf_clk net6 VPWR VGND sg13g2_mux2_1
XFILLER_9_93 VPWR VGND sg13g2_fill_1
X_4665_ net686 net737 _0218_ VPWR VGND sg13g2_nor2_1
X_4755__84 VPWR VGND net84 sg13g2_tiehi
X_4596_ net653 net704 _0149_ VPWR VGND sg13g2_nor2_1
X_3616_ net614 _1340_ _1345_ _1346_ VPWR VGND sg13g2_nor3_1
X_4817__342 VPWR VGND net342 sg13g2_tiehi
X_3547_ net594 VPWR _1277_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\]
+ net586 sg13g2_o21ai_1
X_3478_ _1208_ _1192_ _1196_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_36 VPWR VGND sg13g2_decap_8
X_5079_ net369 VGND VPWR _0626_ tmds_blue.dc_balancing_reg\[3\] net643 sg13g2_dfrbpq_2
XFILLER_44_317 VPWR VGND sg13g2_fill_1
XFILLER_44_306 VPWR VGND sg13g2_decap_4
XFILLER_37_380 VPWR VGND sg13g2_fill_1
XFILLER_25_542 VPWR VGND sg13g2_fill_2
X_4824__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_25_553 VPWR VGND sg13g2_fill_1
XFILLER_13_748 VPWR VGND sg13g2_decap_8
XFILLER_5_925 VPWR VGND sg13g2_decap_8
X_4831__328 VPWR VGND net328 sg13g2_tiehi
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_48_634 VPWR VGND sg13g2_decap_8
XFILLER_47_199 VPWR VGND sg13g2_decap_4
XFILLER_35_339 VPWR VGND sg13g2_decap_4
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
X_2780_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\] _0756_ _0466_
+ VPWR VGND sg13g2_mux2_1
X_4450_ _2132_ _1991_ _2138_ _2139_ VPWR VGND sg13g2_a21o_1
X_3401_ _1088_ net542 _1125_ _1131_ VPWR VGND sg13g2_nor3_1
X_4381_ tmds_blue.dc_balancing_reg\[1\] tmds_blue.n193 _2073_ VPWR VGND sg13g2_xor2_1
X_3332_ _1050_ VPWR _1062_ VGND _1049_ _1051_ sg13g2_o21ai_1
X_4752__87 VPWR VGND net87 sg13g2_tiehi
Xfanout709 net711 net709 VPWR VGND sg13g2_buf_2
X_3263_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ _0367_ _0996_ sg13g2_a21oi_1
X_5002_ net187 VGND VPWR _0549_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\]
+ _0197_ sg13g2_dfrbpq_1
X_3194_ _0802_ _0951_ _0952_ _0334_ VPWR VGND sg13g2_nor3_1
XFILLER_22_1005 VPWR VGND sg13g2_decap_8
XFILLER_38_122 VPWR VGND sg13g2_fill_2
XFILLER_41_309 VPWR VGND sg13g2_decap_8
XFILLER_35_895 VPWR VGND sg13g2_decap_4
X_2978_ VGND VPWR _0818_ _0824_ net17 _0820_ sg13g2_a21oi_1
X_4717_ net149 VGND VPWR _0268_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\]
+ _0007_ sg13g2_dfrbpq_1
X_4648_ net670 net721 _0201_ VPWR VGND sg13g2_nor2_1
X_4579_ net663 net714 _0132_ VPWR VGND sg13g2_nor2_1
XFILLER_39_46 VPWR VGND sg13g2_decap_4
XFILLER_39_79 VPWR VGND sg13g2_decap_8
X_4928__112 VPWR VGND net112 sg13g2_tiehi
XFILLER_29_133 VPWR VGND sg13g2_fill_1
X_4898__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_26_884 VPWR VGND sg13g2_decap_8
XFILLER_13_512 VPWR VGND sg13g2_fill_2
XFILLER_9_505 VPWR VGND sg13g2_decap_8
XFILLER_4_232 VPWR VGND sg13g2_fill_2
XFILLER_5_777 VPWR VGND sg13g2_decap_4
XFILLER_1_972 VPWR VGND sg13g2_decap_8
XFILLER_49_932 VPWR VGND sg13g2_decap_8
XFILLER_48_486 VPWR VGND sg13g2_decap_8
XFILLER_35_114 VPWR VGND sg13g2_decap_8
X_3950_ _1629_ _1658_ _1676_ VPWR VGND sg13g2_nor2_1
XFILLER_16_361 VPWR VGND sg13g2_fill_2
X_2901_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\] _0784_ _0299_
+ VPWR VGND sg13g2_mux2_1
X_3881_ net620 VPWR _1610_ VGND _1608_ _1609_ sg13g2_o21ai_1
X_2832_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\] net763 _0769_ _0427_
+ VPWR VGND sg13g2_mux2_1
X_2763_ net756 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\] _0753_ _0480_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_560 VPWR VGND sg13g2_decap_4
X_4502_ net656 net707 _0055_ VPWR VGND sg13g2_nor2_1
X_2694_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\] _0738_ _0543_
+ VPWR VGND sg13g2_mux2_1
XFILLER_6_61 VPWR VGND sg13g2_fill_1
X_4433_ _2123_ _2101_ _2111_ VPWR VGND sg13g2_nand2_1
XFILLER_6_94 VPWR VGND sg13g2_fill_2
X_4364_ _2059_ _2031_ _2058_ VPWR VGND sg13g2_xnor2_1
X_4295_ tmds_blue.dc_balancing_reg\[4\] _1997_ _1998_ VPWR VGND sg13g2_nor2_2
X_3315_ _1045_ _1042_ _1044_ VPWR VGND sg13g2_nand2_1
X_3246_ _0985_ _0986_ _0360_ VPWR VGND sg13g2_nor2_1
XFILLER_39_453 VPWR VGND sg13g2_decap_4
X_3177_ _0942_ _0794_ _0941_ VPWR VGND sg13g2_nand2_1
XFILLER_27_615 VPWR VGND sg13g2_decap_8
X_4821__338 VPWR VGND net338 sg13g2_tiehi
XFILLER_10_559 VPWR VGND sg13g2_decap_8
XFILLER_6_519 VPWR VGND sg13g2_fill_2
XFILLER_2_758 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_fill_2
XFILLER_46_935 VPWR VGND sg13g2_decap_8
XFILLER_45_478 VPWR VGND sg13g2_fill_2
XFILLER_45_467 VPWR VGND sg13g2_decap_8
XFILLER_33_607 VPWR VGND sg13g2_decap_8
XFILLER_33_618 VPWR VGND sg13g2_fill_1
X_5054__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_26_670 VPWR VGND sg13g2_decap_8
XFILLER_32_106 VPWR VGND sg13g2_fill_2
X_5002__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_32_139 VPWR VGND sg13g2_decap_8
XFILLER_41_684 VPWR VGND sg13g2_decap_4
XFILLER_41_662 VPWR VGND sg13g2_decap_4
XFILLER_9_368 VPWR VGND sg13g2_fill_2
XFILLER_31_91 VPWR VGND sg13g2_decap_8
X_3100_ _0890_ _0884_ _0889_ VPWR VGND sg13g2_nand2_1
XFILLER_49_751 VPWR VGND sg13g2_decap_8
X_4080_ VPWR _1803_ _1802_ VGND sg13g2_inv_1
X_5083__248 VPWR VGND net248 sg13g2_tiehi
X_3031_ net419 red_tmds_par\[6\] net696 serialize.n427\[6\] VPWR VGND sg13g2_mux2_1
X_4727__136 VPWR VGND net136 sg13g2_tiehi
X_4982_ net269 VGND VPWR _0529_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\]
+ _0177_ sg13g2_dfrbpq_1
X_3933_ _1630_ net544 _1659_ VPWR VGND sg13g2_xor2_1
X_3864_ net621 VPWR _1593_ VGND _1591_ _1592_ sg13g2_o21ai_1
X_2815_ _0718_ _0762_ _0766_ VPWR VGND sg13g2_nor2_2
XFILLER_20_846 VPWR VGND sg13g2_fill_1
X_3795_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\] net589 _1525_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_891 VPWR VGND sg13g2_fill_1
X_2746_ _0689_ _0723_ _0749_ VPWR VGND sg13g2_nor2_2
X_2677_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\] _0735_ _0557_
+ VPWR VGND sg13g2_mux2_1
X_4416_ _2106_ tmds_blue.n193 _2105_ VPWR VGND sg13g2_nand2_1
X_4347_ _2042_ _0641_ _2027_ VPWR VGND sg13g2_xnor2_1
X_4278_ _0889_ VPWR _1983_ VGND _1970_ _1982_ sg13g2_o21ai_1
X_3229_ net609 _0897_ _0974_ VPWR VGND sg13g2_and2_1
XFILLER_28_935 VPWR VGND sg13g2_decap_8
XFILLER_27_412 VPWR VGND sg13g2_fill_1
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_43_949 VPWR VGND sg13g2_decap_8
XFILLER_42_437 VPWR VGND sg13g2_fill_1
XFILLER_42_426 VPWR VGND sg13g2_decap_4
XFILLER_14_106 VPWR VGND sg13g2_decap_4
XFILLER_10_301 VPWR VGND sg13g2_decap_8
XFILLER_35_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_389 VPWR VGND sg13g2_decap_4
XFILLER_18_401 VPWR VGND sg13g2_decap_8
XFILLER_19_935 VPWR VGND sg13g2_decap_8
XFILLER_46_765 VPWR VGND sg13g2_fill_1
XFILLER_42_993 VPWR VGND sg13g2_decap_8
X_4804__366 VPWR VGND net366 sg13g2_tiehi
XFILLER_14_684 VPWR VGND sg13g2_fill_2
XFILLER_9_143 VPWR VGND sg13g2_fill_1
XFILLER_9_132 VPWR VGND sg13g2_fill_1
XFILLER_9_121 VPWR VGND sg13g2_decap_8
XFILLER_9_154 VPWR VGND sg13g2_decap_4
X_2600_ VPWR _0707_ _0706_ VGND sg13g2_inv_1
X_3580_ net594 VPWR _1310_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\]
+ net565 sg13g2_o21ai_1
XFILLER_9_187 VPWR VGND sg13g2_decap_8
X_4943__57 VPWR VGND net57 sg13g2_tiehi
X_2531_ _0649_ net600 VPWR VGND sg13g2_inv_8
X_4201_ _1917_ _0889_ _1916_ VPWR VGND sg13g2_xnor2_1
X_4132_ _1850_ _1842_ _1855_ VPWR VGND _1853_ sg13g2_nand3b_1
XFILLER_3_1002 VPWR VGND sg13g2_decap_8
X_4063_ VGND VPWR _1783_ _1785_ _1786_ _1779_ sg13g2_a21oi_1
XFILLER_49_581 VPWR VGND sg13g2_decap_8
X_3014_ net425 green_tmds_par\[0\] net698 serialize.n428\[0\] VPWR VGND sg13g2_mux2_1
XFILLER_25_927 VPWR VGND sg13g2_decap_8
X_4965_ net359 VGND VPWR _0512_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\]
+ _0160_ sg13g2_dfrbpq_1
X_3916_ _1642_ _1084_ _1632_ VPWR VGND sg13g2_nand2_1
X_4740__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_33_993 VPWR VGND sg13g2_decap_8
X_4896_ net204 VGND VPWR _0447_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\]
+ _0104_ sg13g2_dfrbpq_1
X_3847_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\] net590 _1576_ VPWR
+ VGND sg13g2_nor2_1
X_3778_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\] net581 _1508_ VPWR
+ VGND sg13g2_nor2_1
X_2729_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\] net780 _0745_ _0515_
+ VPWR VGND sg13g2_mux2_1
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_15_404 VPWR VGND sg13g2_fill_2
XFILLER_15_415 VPWR VGND sg13g2_fill_2
XFILLER_42_278 VPWR VGND sg13g2_decap_4
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_23_481 VPWR VGND sg13g2_decap_8
XFILLER_23_492 VPWR VGND sg13g2_fill_2
XFILLER_11_654 VPWR VGND sg13g2_decap_4
XFILLER_10_175 VPWR VGND sg13g2_fill_2
XFILLER_7_658 VPWR VGND sg13g2_decap_8
XFILLER_6_113 VPWR VGND sg13g2_decap_4
XFILLER_3_897 VPWR VGND sg13g2_decap_8
XFILLER_38_507 VPWR VGND sg13g2_fill_2
XFILLER_34_724 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_decap_4
X_4724__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_30_930 VPWR VGND sg13g2_decap_8
X_4750_ net91 VGND VPWR _0301_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\]
+ _0032_ sg13g2_dfrbpq_1
X_3701_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\] net553 _1431_ VPWR
+ VGND sg13g2_nor2_1
X_4681_ net663 net714 _0234_ VPWR VGND sg13g2_nor2_1
X_3632_ _1358_ _1359_ _1360_ _1361_ _1362_ VPWR VGND sg13g2_nor4_1
X_3563_ net594 VPWR _1293_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\]
+ net566 sg13g2_o21ai_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2514_ VPWR _0632_ videogen.fancy_shader.video_y\[9\] VGND sg13g2_inv_1
X_3494_ _1212_ _1204_ _1224_ VPWR VGND _1222_ sg13g2_nand3b_1
XFILLER_25_1025 VPWR VGND sg13g2_decap_4
X_4115_ _1838_ _1802_ _1837_ VPWR VGND sg13g2_nand2_1
X_5095_ net801 VGND VPWR serialize.n431\[0\] serialize.n459 clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_2537__1 VPWR net405 clknet_1_0__leaf_clk VGND sg13g2_inv_1
X_4046_ _1769_ _1728_ _1766_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_16 VPWR VGND sg13g2_decap_8
XFILLER_37_584 VPWR VGND sg13g2_fill_2
XFILLER_24_223 VPWR VGND sg13g2_decap_4
XFILLER_12_418 VPWR VGND sg13g2_fill_1
X_4948_ net37 VGND VPWR _0495_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\]
+ _0152_ sg13g2_dfrbpq_1
X_4879_ net237 VGND VPWR _0430_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\]
+ _0087_ sg13g2_dfrbpq_1
XFILLER_32_1018 VPWR VGND sg13g2_decap_8
XFILLER_21_985 VPWR VGND sg13g2_decap_8
XFILLER_0_856 VPWR VGND sg13g2_decap_8
XFILLER_28_562 VPWR VGND sg13g2_fill_1
XFILLER_15_245 VPWR VGND sg13g2_fill_1
XFILLER_15_267 VPWR VGND sg13g2_decap_4
XFILLER_8_912 VPWR VGND sg13g2_decap_8
XFILLER_12_974 VPWR VGND sg13g2_decap_8
X_4749__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_8_989 VPWR VGND sg13g2_decap_8
XFILLER_48_1014 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_fill_1
XFILLER_38_359 VPWR VGND sg13g2_fill_1
XFILLER_38_348 VPWR VGND sg13g2_fill_1
XFILLER_19_551 VPWR VGND sg13g2_decap_8
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_85 VPWR VGND sg13g2_decap_4
XFILLER_19_595 VPWR VGND sg13g2_decap_4
X_2994_ serialize.n455 serialize.n453 clknet_1_1__leaf_clk net5 VPWR VGND sg13g2_mux2_1
X_4802_ net370 VGND VPWR _0353_ videogen.fancy_shader.n646\[7\] net633 sg13g2_dfrbpq_2
XFILLER_9_50 VPWR VGND sg13g2_decap_8
X_4733_ net125 VGND VPWR _0284_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\]
+ _0015_ sg13g2_dfrbpq_1
X_4664_ net676 net728 _0217_ VPWR VGND sg13g2_nor2_1
X_4595_ net655 net706 _0148_ VPWR VGND sg13g2_nor2_1
X_3615_ _1341_ _1342_ _1343_ _1344_ _1345_ VPWR VGND sg13g2_nor4_1
X_3546_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] VPWR _1276_ VGND _1269_
+ _1275_ sg13g2_o21ai_1
X_3477_ _1195_ _1201_ _1056_ _1207_ VPWR VGND _1202_ sg13g2_nand4_1
XFILLER_29_315 VPWR VGND sg13g2_fill_1
X_5078_ net31 VGND VPWR _0625_ tmds_blue.dc_balancing_reg\[2\] net641 sg13g2_dfrbpq_1
X_4029_ _1752_ _1633_ _1751_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_524 VPWR VGND sg13g2_decap_8
XFILLER_12_204 VPWR VGND sg13g2_fill_1
XFILLER_12_226 VPWR VGND sg13g2_fill_1
XFILLER_13_727 VPWR VGND sg13g2_decap_4
XFILLER_25_598 VPWR VGND sg13g2_decap_8
XFILLER_12_259 VPWR VGND sg13g2_fill_1
XFILLER_5_904 VPWR VGND sg13g2_decap_8
XFILLER_21_793 VPWR VGND sg13g2_decap_8
XFILLER_5_19 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_30 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_0_642 VPWR VGND sg13g2_decap_8
X_4868__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_47_189 VPWR VGND sg13g2_fill_1
XFILLER_18_70 VPWR VGND sg13g2_decap_8
XFILLER_28_381 VPWR VGND sg13g2_decap_8
XFILLER_7_241 VPWR VGND sg13g2_decap_4
X_4875__245 VPWR VGND net245 sg13g2_tiehi
XFILLER_12_793 VPWR VGND sg13g2_decap_8
X_3400_ VGND VPWR _1115_ _1120_ _1130_ _1124_ sg13g2_a21oi_1
X_4380_ net749 clockdiv.q0 net406 _0623_ VPWR VGND sg13g2_nor3_1
X_3331_ _1061_ videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.n646\[5\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_4_992 VPWR VGND sg13g2_decap_8
XFILLER_39_602 VPWR VGND sg13g2_fill_1
X_3262_ net793 VPWR _0996_ VGND videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ sg13g2_o21ai_1
X_3193_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0792_ _0952_ VPWR
+ VGND sg13g2_nor2_1
X_4847__303 VPWR VGND net303 sg13g2_tiehi
X_5001_ net191 VGND VPWR _0548_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\]
+ _0196_ sg13g2_dfrbpq_1
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_38_156 VPWR VGND sg13g2_fill_1
XFILLER_26_318 VPWR VGND sg13g2_fill_1
XFILLER_14_39 VPWR VGND sg13g2_fill_1
X_2977_ _0824_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0822_ VPWR VGND
+ sg13g2_xnor2_1
X_4716_ net151 VGND VPWR _0267_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\]
+ _0006_ sg13g2_dfrbpq_1
X_4647_ net668 net720 _0200_ VPWR VGND sg13g2_nor2_1
X_4578_ net664 net715 _0131_ VPWR VGND sg13g2_nor2_1
X_3529_ net594 VPWR _1259_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\]
+ net577 sg13g2_o21ai_1
XFILLER_29_101 VPWR VGND sg13g2_fill_1
XFILLER_44_159 VPWR VGND sg13g2_decap_8
XFILLER_25_351 VPWR VGND sg13g2_decap_8
XFILLER_40_310 VPWR VGND sg13g2_decap_8
XFILLER_41_855 VPWR VGND sg13g2_fill_2
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_5_756 VPWR VGND sg13g2_decap_4
XFILLER_45_1006 VPWR VGND sg13g2_decap_8
XFILLER_4_299 VPWR VGND sg13g2_decap_4
XFILLER_1_951 VPWR VGND sg13g2_decap_8
XFILLER_49_911 VPWR VGND sg13g2_decap_8
XFILLER_0_450 VPWR VGND sg13g2_fill_1
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_49_988 VPWR VGND sg13g2_decap_8
XFILLER_17_841 VPWR VGND sg13g2_fill_2
X_2900_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\] _0784_ _0300_
+ VPWR VGND sg13g2_mux2_1
X_3880_ _1564_ VPWR _1609_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\]
+ net585 sg13g2_o21ai_1
X_2831_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\] net753 _0769_ _0428_
+ VPWR VGND sg13g2_mux2_1
X_2762_ _0753_ _0710_ _0751_ VPWR VGND sg13g2_nand2_2
X_4501_ net651 net702 _0054_ VPWR VGND sg13g2_nor2_1
X_4432_ _2122_ _2097_ _2119_ VPWR VGND sg13g2_xnor2_1
X_2693_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\] _0738_ _0544_
+ VPWR VGND sg13g2_mux2_1
X_4814__346 VPWR VGND net346 sg13g2_tiehi
X_4363_ _2058_ _2042_ _2056_ VPWR VGND sg13g2_xnor2_1
X_4294_ net606 VPWR _1997_ VGND _1988_ _1996_ sg13g2_o21ai_1
X_3314_ videogen.fancy_shader.video_x\[4\] videogen.fancy_shader.n646\[4\] _1044_
+ VPWR VGND sg13g2_xor2_1
X_3245_ net795 VPWR _0986_ VGND videogen.fancy_shader.video_y\[4\] _0984_ sg13g2_o21ai_1
X_3176_ net616 _0938_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] _0941_
+ VPWR VGND sg13g2_nand3_1
XFILLER_27_638 VPWR VGND sg13g2_decap_4
XFILLER_23_833 VPWR VGND sg13g2_decap_8
XFILLER_35_682 VPWR VGND sg13g2_fill_1
XFILLER_23_899 VPWR VGND sg13g2_decap_8
XFILLER_41_37 VPWR VGND sg13g2_decap_8
XFILLER_46_914 VPWR VGND sg13g2_decap_8
XFILLER_18_616 VPWR VGND sg13g2_decap_8
XFILLER_45_435 VPWR VGND sg13g2_fill_1
XFILLER_17_159 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_fill_2
XFILLER_13_398 VPWR VGND sg13g2_decap_8
XFILLER_12_1016 VPWR VGND sg13g2_decap_8
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_5_597 VPWR VGND sg13g2_fill_1
XFILLER_49_730 VPWR VGND sg13g2_decap_8
XFILLER_0_291 VPWR VGND sg13g2_decap_4
X_3030_ net423 red_tmds_par\[5\] net697 serialize.n427\[5\] VPWR VGND sg13g2_mux2_1
X_4981_ net273 VGND VPWR _0528_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\]
+ _0176_ sg13g2_dfrbpq_1
XFILLER_17_682 VPWR VGND sg13g2_decap_8
X_3932_ _1658_ _1635_ _1656_ VPWR VGND sg13g2_xnor2_1
X_3863_ _1570_ VPWR _1592_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\]
+ net587 sg13g2_o21ai_1
XFILLER_31_151 VPWR VGND sg13g2_decap_8
X_2814_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\] net785 _0765_ _0441_
+ VPWR VGND sg13g2_mux2_1
X_3794_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\] net580 _1524_ VPWR
+ VGND sg13g2_nor2_1
X_2745_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\] _0748_ _0493_
+ VPWR VGND sg13g2_mux2_1
X_2676_ _0735_ _0702_ _0731_ VPWR VGND sg13g2_nand2_2
X_4415_ _2105_ net604 _2077_ VPWR VGND sg13g2_nand2_1
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
X_4346_ _2018_ _2029_ _2041_ VPWR VGND sg13g2_nor2_1
X_4277_ _1982_ _1979_ _1981_ VPWR VGND sg13g2_xnor2_1
X_3228_ net747 _0972_ _0973_ _0355_ VPWR VGND sg13g2_nor3_1
XFILLER_28_914 VPWR VGND sg13g2_decap_8
X_3159_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\] _0928_ _0929_
+ _0919_ sg13g2_a21oi_1
XFILLER_27_435 VPWR VGND sg13g2_decap_4
XFILLER_43_928 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_35_1005 VPWR VGND sg13g2_decap_8
XFILLER_11_847 VPWR VGND sg13g2_decap_4
XFILLER_2_578 VPWR VGND sg13g2_decap_4
XFILLER_18_446 VPWR VGND sg13g2_fill_2
XFILLER_34_928 VPWR VGND sg13g2_fill_1
XFILLER_42_972 VPWR VGND sg13g2_decap_8
X_2530_ _0648_ net793 VPWR VGND sg13g2_inv_2
X_4200_ _1916_ tmds_red.n126 _0860_ VPWR VGND sg13g2_xnor2_1
X_4131_ _1843_ VPWR _1854_ VGND _1851_ _1853_ sg13g2_o21ai_1
XFILLER_49_560 VPWR VGND sg13g2_decap_8
X_4062_ _1785_ _1774_ _1784_ VPWR VGND sg13g2_nand2_1
X_3013_ blue_tmds_par\[9\] net696 serialize.n429\[9\] VPWR VGND sg13g2_and2_1
XFILLER_37_733 VPWR VGND sg13g2_decap_4
XFILLER_37_755 VPWR VGND sg13g2_fill_1
XFILLER_25_906 VPWR VGND sg13g2_decap_8
XFILLER_18_980 VPWR VGND sg13g2_decap_8
X_4964_ net363 VGND VPWR _0511_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\]
+ _0159_ sg13g2_dfrbpq_1
X_3915_ _1641_ _1087_ _1632_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_972 VPWR VGND sg13g2_decap_8
X_4895_ net206 VGND VPWR _0446_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\]
+ _0103_ sg13g2_dfrbpq_1
X_3846_ _1574_ VPWR _1575_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\]
+ net589 sg13g2_o21ai_1
X_3777_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\] net587 _1507_ VPWR
+ VGND sg13g2_nor2_1
X_2728_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\] net769 _0745_ _0516_
+ VPWR VGND sg13g2_mux2_1
X_2659_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\] _0730_ _0570_
+ VPWR VGND sg13g2_mux2_1
X_4329_ net602 _2021_ _2025_ VPWR VGND sg13g2_nor2_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_755 VPWR VGND sg13g2_fill_1
XFILLER_43_703 VPWR VGND sg13g2_fill_1
XFILLER_42_224 VPWR VGND sg13g2_fill_2
XFILLER_15_449 VPWR VGND sg13g2_decap_8
XFILLER_30_419 VPWR VGND sg13g2_fill_1
X_4776__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_11_666 VPWR VGND sg13g2_fill_1
XFILLER_10_187 VPWR VGND sg13g2_decap_8
XFILLER_10_198 VPWR VGND sg13g2_fill_1
XFILLER_3_821 VPWR VGND sg13g2_decap_8
XFILLER_3_876 VPWR VGND sg13g2_decap_8
Xfanout690 net691 net690 VPWR VGND sg13g2_buf_8
XFILLER_18_221 VPWR VGND sg13g2_fill_1
XFILLER_37_80 VPWR VGND sg13g2_decap_8
XFILLER_18_276 VPWR VGND sg13g2_fill_2
XFILLER_19_788 VPWR VGND sg13g2_decap_8
XFILLER_34_703 VPWR VGND sg13g2_decap_8
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
XFILLER_14_460 VPWR VGND sg13g2_decap_8
XFILLER_15_994 VPWR VGND sg13g2_decap_8
X_3700_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\] net563 _1430_ VPWR
+ VGND sg13g2_nor2_1
X_4680_ net671 net722 _0233_ VPWR VGND sg13g2_nor2_1
XFILLER_30_986 VPWR VGND sg13g2_decap_8
X_3631_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\] net565 _1361_ VPWR
+ VGND sg13g2_nor2_1
X_3562_ _1288_ _1289_ _1290_ _1291_ _1292_ VPWR VGND sg13g2_nor4_1
X_3493_ _1203_ VPWR _1223_ VGND _1213_ _1222_ sg13g2_o21ai_1
X_4989__238 VPWR VGND net238 sg13g2_tiehi
XFILLER_38_0 VPWR VGND sg13g2_decap_4
XFILLER_25_1004 VPWR VGND sg13g2_decap_8
X_4114_ _1835_ _1832_ _1836_ _1837_ VPWR VGND sg13g2_a21o_2
X_5094_ net801 VGND VPWR serialize.n428\[9\] serialize.n414\[7\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4045_ _1766_ _1728_ _1768_ VPWR VGND sg13g2_xor2_1
XFILLER_24_202 VPWR VGND sg13g2_decap_8
XFILLER_12_408 VPWR VGND sg13g2_fill_1
X_4947_ net41 VGND VPWR _0494_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\]
+ _0151_ sg13g2_dfrbpq_1
X_4878_ net239 VGND VPWR _0429_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\]
+ _0086_ sg13g2_dfrbpq_1
XFILLER_21_964 VPWR VGND sg13g2_decap_8
X_3829_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\] net588 _1558_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_474 VPWR VGND sg13g2_decap_8
XFILLER_3_117 VPWR VGND sg13g2_fill_1
XFILLER_0_835 VPWR VGND sg13g2_decap_8
XFILLER_48_828 VPWR VGND sg13g2_fill_2
XFILLER_16_714 VPWR VGND sg13g2_decap_8
XFILLER_28_552 VPWR VGND sg13g2_fill_1
XFILLER_16_758 VPWR VGND sg13g2_decap_8
XFILLER_24_791 VPWR VGND sg13g2_fill_2
X_4723__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_12_953 VPWR VGND sg13g2_decap_8
XFILLER_11_452 VPWR VGND sg13g2_decap_4
XFILLER_8_968 VPWR VGND sg13g2_decap_8
XFILLER_3_640 VPWR VGND sg13g2_decap_8
XFILLER_3_651 VPWR VGND sg13g2_fill_1
XFILLER_3_684 VPWR VGND sg13g2_decap_8
XFILLER_38_327 VPWR VGND sg13g2_fill_1
XFILLER_0_53 VPWR VGND sg13g2_fill_2
XFILLER_0_1017 VPWR VGND sg13g2_decap_8
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
XFILLER_34_544 VPWR VGND sg13g2_decap_4
XFILLER_34_566 VPWR VGND sg13g2_fill_2
X_2993_ serialize.n458 serialize.n456 clknet_1_0__leaf_clk net3 VPWR VGND sg13g2_mux2_1
X_4801_ net372 VGND VPWR _0352_ videogen.fancy_shader.n646\[6\] net638 sg13g2_dfrbpq_2
XFILLER_21_205 VPWR VGND sg13g2_decap_8
X_4732_ net127 VGND VPWR _0283_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\]
+ _0014_ sg13g2_dfrbpq_1
X_4663_ net659 net710 _0216_ VPWR VGND sg13g2_nor2_1
X_3614_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\] net584 _1344_ VPWR
+ VGND sg13g2_nor2_1
X_4594_ net655 net706 _0147_ VPWR VGND sg13g2_nor2_1
X_3545_ net614 VPWR _1275_ VGND _1270_ _1274_ sg13g2_o21ai_1
X_3476_ _1206_ _1195_ _1201_ VPWR VGND sg13g2_xnor2_1
X_5063__225 VPWR VGND net225 sg13g2_tiehi
X_5077_ net47 VGND VPWR _0624_ tmds_blue.dc_balancing_reg\[1\] net641 sg13g2_dfrbpq_2
X_4028_ VGND VPWR _1060_ _1750_ _1751_ _1729_ sg13g2_a21oi_1
XFILLER_25_511 VPWR VGND sg13g2_fill_1
XFILLER_12_238 VPWR VGND sg13g2_fill_1
XFILLER_4_404 VPWR VGND sg13g2_fill_1
X_4761__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_0_632 VPWR VGND sg13g2_fill_2
XFILLER_48_625 VPWR VGND sg13g2_decap_4
X_5081__314 VPWR VGND net314 sg13g2_tiehi
XFILLER_47_135 VPWR VGND sg13g2_fill_2
XFILLER_29_850 VPWR VGND sg13g2_fill_1
XFILLER_47_168 VPWR VGND sg13g2_decap_8
X_5005__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_12_761 VPWR VGND sg13g2_fill_1
XFILLER_4_971 VPWR VGND sg13g2_decap_8
X_3330_ _1060_ _1058_ _1059_ VPWR VGND sg13g2_xnor2_1
X_5000_ net195 VGND VPWR _0547_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\]
+ _0195_ sg13g2_dfrbpq_1
X_3261_ videogen.test_lut_thingy.gol_counter_reg\[0\] net749 _0366_ VPWR VGND sg13g2_nor2_1
X_3192_ _0794_ VPWR _0951_ VGND _0931_ _0932_ sg13g2_o21ai_1
XFILLER_38_124 VPWR VGND sg13g2_fill_1
XFILLER_22_569 VPWR VGND sg13g2_decap_8
X_2976_ VGND VPWR _0818_ _0823_ net16 _0820_ sg13g2_a21oi_1
X_4715_ net152 VGND VPWR net737 clockdiv.q2temp net405 sg13g2_dfrbpq_1
X_4646_ net670 net721 _0199_ VPWR VGND sg13g2_nor2_1
X_4737__117 VPWR VGND net117 sg13g2_tiehi
X_4577_ net661 net712 _0130_ VPWR VGND sg13g2_nor2_1
X_3528_ _1252_ _1254_ _1256_ _1257_ _1258_ VPWR VGND sg13g2_nor4_1
X_3459_ _1184_ _1185_ _1180_ _1189_ VPWR VGND sg13g2_nand3_1
XFILLER_18_809 VPWR VGND sg13g2_fill_2
XFILLER_29_113 VPWR VGND sg13g2_fill_2
XFILLER_38_1014 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
X_4720__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_40_366 VPWR VGND sg13g2_decap_4
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_4_278 VPWR VGND sg13g2_decap_8
XFILLER_1_930 VPWR VGND sg13g2_decap_8
XFILLER_48_400 VPWR VGND sg13g2_decap_8
XFILLER_49_967 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_fill_1
XFILLER_29_92 VPWR VGND sg13g2_fill_2
XFILLER_17_820 VPWR VGND sg13g2_fill_2
XFILLER_16_330 VPWR VGND sg13g2_fill_2
XFILLER_28_190 VPWR VGND sg13g2_fill_1
XFILLER_45_80 VPWR VGND sg13g2_decap_8
X_2830_ _0725_ _0762_ _0769_ VPWR VGND sg13g2_nor2_2
XFILLER_31_333 VPWR VGND sg13g2_fill_2
XFILLER_32_867 VPWR VGND sg13g2_decap_4
X_2761_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\] _0752_ _0481_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_388 VPWR VGND sg13g2_decap_8
XFILLER_31_399 VPWR VGND sg13g2_fill_2
X_2692_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\] _0738_ _0545_
+ VPWR VGND sg13g2_mux2_1
X_4500_ net652 net703 _0053_ VPWR VGND sg13g2_nor2_1
X_4957__387 VPWR VGND net387 sg13g2_tiehi
X_4431_ VGND VPWR _2004_ _2113_ _2121_ _2120_ sg13g2_a21oi_1
X_4362_ _2043_ _2056_ _2057_ VPWR VGND sg13g2_nor2_1
X_3313_ _1043_ videogen.fancy_shader.n646\[4\] videogen.fancy_shader.video_x\[4\]
+ VPWR VGND sg13g2_nand2_1
X_4293_ _1996_ net604 tmds_blue.n193 VPWR VGND sg13g2_xnor2_1
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
X_3244_ _0816_ _0976_ _0985_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_1023 VPWR VGND sg13g2_fill_2
XFILLER_20_0 VPWR VGND sg13g2_fill_1
X_3175_ VGND VPWR net616 _0938_ _0940_ net613 sg13g2_a21oi_1
XFILLER_23_812 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_23_878 VPWR VGND sg13g2_decap_8
X_2959_ VGND VPWR _0649_ net8 _0671_ net627 sg13g2_a21oi_2
XFILLER_22_388 VPWR VGND sg13g2_fill_2
X_4629_ net689 net741 _0182_ VPWR VGND sg13g2_nor2_1
XFILLER_2_727 VPWR VGND sg13g2_fill_1
XFILLER_2_716 VPWR VGND sg13g2_decap_8
XFILLER_1_237 VPWR VGND sg13g2_fill_2
XFILLER_26_650 VPWR VGND sg13g2_fill_2
XFILLER_26_694 VPWR VGND sg13g2_fill_2
XFILLER_13_366 VPWR VGND sg13g2_fill_1
XFILLER_40_196 VPWR VGND sg13g2_fill_2
XFILLER_5_554 VPWR VGND sg13g2_fill_2
Xoutput3 net3 tmds_b VPWR VGND sg13g2_buf_1
XFILLER_0_270 VPWR VGND sg13g2_decap_8
XFILLER_36_414 VPWR VGND sg13g2_decap_4
XFILLER_36_469 VPWR VGND sg13g2_decap_8
XFILLER_45_992 VPWR VGND sg13g2_decap_8
XFILLER_23_119 VPWR VGND sg13g2_decap_8
X_4980_ net277 VGND VPWR _0527_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\]
+ _0175_ sg13g2_dfrbpq_1
X_3931_ _1657_ _1634_ _1656_ VPWR VGND sg13g2_xnor2_1
X_3862_ _1569_ VPWR _1591_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\]
+ net578 sg13g2_o21ai_1
XFILLER_32_675 VPWR VGND sg13g2_decap_4
X_2813_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\] net773 _0765_ _0442_
+ VPWR VGND sg13g2_mux2_1
X_4946__45 VPWR VGND net45 sg13g2_tiehi
X_3793_ net597 VPWR _1523_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\]
+ net566 sg13g2_o21ai_1
XFILLER_9_882 VPWR VGND sg13g2_decap_8
X_2744_ net772 videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\] _0748_ _0494_
+ VPWR VGND sg13g2_mux2_1
X_2675_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\] _0734_ _0558_
+ VPWR VGND sg13g2_mux2_1
X_4414_ _2085_ _2087_ _2104_ VPWR VGND sg13g2_nor2_1
X_4345_ net569 _2040_ _0620_ VPWR VGND sg13g2_nor2_1
X_4276_ _1981_ tmds_red.dc_balancing_reg\[4\] _1980_ VPWR VGND sg13g2_xnor2_1
X_3227_ _0973_ videogen.fancy_shader.n646\[9\] videogen.fancy_shader.n646\[8\] _0970_
+ VPWR VGND sg13g2_and3_1
XFILLER_39_285 VPWR VGND sg13g2_decap_4
XFILLER_39_274 VPWR VGND sg13g2_decap_8
X_3158_ _0919_ _0927_ _0928_ _0322_ VPWR VGND sg13g2_nor3_1
XFILLER_43_907 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
X_3089_ _0879_ _0877_ _0876_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_970 VPWR VGND sg13g2_fill_1
XFILLER_22_130 VPWR VGND sg13g2_fill_1
XFILLER_35_1028 VPWR VGND sg13g2_fill_1
XFILLER_23_697 VPWR VGND sg13g2_fill_2
XFILLER_7_819 VPWR VGND sg13g2_decap_8
XFILLER_10_336 VPWR VGND sg13g2_decap_8
X_4901__194 VPWR VGND net194 sg13g2_tiehi
X_5036__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_7_4 VPWR VGND sg13g2_fill_2
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_2_568 VPWR VGND sg13g2_fill_2
X_5082__283 VPWR VGND net283 sg13g2_tiehi
XFILLER_46_789 VPWR VGND sg13g2_decap_8
XFILLER_26_82 VPWR VGND sg13g2_decap_8
XFILLER_33_439 VPWR VGND sg13g2_fill_2
XFILLER_42_951 VPWR VGND sg13g2_decap_8
XFILLER_14_686 VPWR VGND sg13g2_fill_1
XFILLER_10_881 VPWR VGND sg13g2_fill_1
XFILLER_6_863 VPWR VGND sg13g2_decap_4
XFILLER_5_340 VPWR VGND sg13g2_decap_8
X_4130_ VGND VPWR _1832_ _1835_ _1853_ _1852_ sg13g2_a21oi_1
XFILLER_3_20 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_3_97 VPWR VGND sg13g2_decap_8
X_4061_ _1781_ VPWR _1784_ VGND _1769_ _1777_ sg13g2_o21ai_1
X_3012_ blue_tmds_par\[8\] net695 serialize.n429\[8\] VPWR VGND sg13g2_and2_1
XFILLER_36_244 VPWR VGND sg13g2_decap_8
X_4963_ net367 VGND VPWR _0510_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\]
+ _0158_ sg13g2_dfrbpq_1
X_3914_ _1640_ net542 _1638_ VPWR VGND sg13g2_xnor2_1
X_4894_ net208 VGND VPWR _0445_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\]
+ _0102_ sg13g2_dfrbpq_1
XFILLER_20_612 VPWR VGND sg13g2_fill_2
X_3845_ _1572_ _1573_ _1574_ VPWR VGND sg13g2_nor2_1
X_3776_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\] net563 _1506_ VPWR
+ VGND sg13g2_nor2_1
X_2727_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\] net759 _0745_ _0517_
+ VPWR VGND sg13g2_mux2_1
X_4855__288 VPWR VGND net288 sg13g2_tiehi
X_2658_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\] _0730_ _0571_
+ VPWR VGND sg13g2_mux2_1
X_5066__201 VPWR VGND net201 sg13g2_tiehi
X_2589_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\] net782 _0700_ _0628_
+ VPWR VGND sg13g2_mux2_1
X_4328_ tmds_green.n132 tmds_green.n126 net603 _2024_ VPWR VGND sg13g2_nand3_1
XFILLER_41_1021 VPWR VGND sg13g2_decap_8
X_4259_ _1965_ _1955_ _1964_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_723 VPWR VGND sg13g2_decap_4
XFILLER_27_233 VPWR VGND sg13g2_fill_2
XFILLER_16_929 VPWR VGND sg13g2_decap_8
XFILLER_27_266 VPWR VGND sg13g2_fill_1
XFILLER_15_428 VPWR VGND sg13g2_decap_8
XFILLER_11_623 VPWR VGND sg13g2_fill_2
XFILLER_24_995 VPWR VGND sg13g2_decap_8
Xfanout691 net692 net691 VPWR VGND sg13g2_buf_8
Xfanout680 net683 net680 VPWR VGND sg13g2_buf_8
XFILLER_19_712 VPWR VGND sg13g2_decap_8
XFILLER_19_756 VPWR VGND sg13g2_decap_8
XFILLER_19_767 VPWR VGND sg13g2_fill_1
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_33_258 VPWR VGND sg13g2_fill_1
XFILLER_30_965 VPWR VGND sg13g2_decap_8
X_3630_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\] net588 _1360_ VPWR
+ VGND sg13g2_nor2_1
X_3561_ net622 VPWR _1291_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\]
+ net580 sg13g2_o21ai_1
X_3492_ VPWR VGND _1216_ _1215_ _1211_ _1034_ _1222_ _1035_ sg13g2_a221oi_1
X_5093_ net798 VGND VPWR serialize.n428\[8\] serialize.n414\[6\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4113_ _1828_ _1823_ _1827_ _1836_ VPWR VGND sg13g2_mux2_1
X_4885__226 VPWR VGND net226 sg13g2_tiehi
XFILLER_29_509 VPWR VGND sg13g2_fill_2
XFILLER_49_380 VPWR VGND sg13g2_decap_8
XFILLER_37_531 VPWR VGND sg13g2_decap_8
X_4044_ _1728_ _1766_ _1767_ VPWR VGND sg13g2_nor2_1
XFILLER_37_597 VPWR VGND sg13g2_fill_2
XFILLER_37_586 VPWR VGND sg13g2_fill_1
XFILLER_25_748 VPWR VGND sg13g2_fill_2
X_4946_ net45 VGND VPWR _0493_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\]
+ _0150_ sg13g2_dfrbpq_1
X_4877_ net241 VGND VPWR _0428_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\]
+ _0085_ sg13g2_dfrbpq_1
XFILLER_21_943 VPWR VGND sg13g2_decap_8
X_3828_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\] net555 _1557_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_453 VPWR VGND sg13g2_fill_2
XFILLER_20_497 VPWR VGND sg13g2_decap_4
X_3759_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\] net552 _1489_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_814 VPWR VGND sg13g2_decap_8
XFILLER_28_531 VPWR VGND sg13g2_fill_1
XFILLER_43_534 VPWR VGND sg13g2_decap_8
XFILLER_28_597 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_fill_2
XFILLER_15_236 VPWR VGND sg13g2_fill_1
XFILLER_12_932 VPWR VGND sg13g2_decap_8
XFILLER_8_947 VPWR VGND sg13g2_decap_8
XFILLER_11_497 VPWR VGND sg13g2_fill_2
XFILLER_3_663 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_34_501 VPWR VGND sg13g2_fill_1
X_4800_ net374 VGND VPWR _0351_ videogen.fancy_shader.n646\[5\] net636 sg13g2_dfrbpq_2
X_2992_ serialize.n461 serialize.n459 clknet_1_0__leaf_clk net4 VPWR VGND sg13g2_mux2_1
XFILLER_22_729 VPWR VGND sg13g2_decap_4
XFILLER_34_578 VPWR VGND sg13g2_decap_8
X_4731_ net129 VGND VPWR _0282_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[3\]
+ _0013_ sg13g2_dfrbpq_1
X_4662_ net659 net710 _0215_ VPWR VGND sg13g2_nor2_1
X_3613_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\] net561 _1343_ VPWR
+ VGND sg13g2_nor2_1
X_4593_ net654 net705 _0146_ VPWR VGND sg13g2_nor2_1
X_3544_ _1273_ VPWR _1274_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[2\]
+ net582 sg13g2_o21ai_1
X_3475_ VPWR VGND _1200_ _1194_ _1197_ _1064_ _1205_ _1065_ sg13g2_a221oi_1
X_4787__400 VPWR VGND net400 sg13g2_tiehi
X_5076_ net63 VGND VPWR net407 clockdiv.q0 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
X_4027_ _1750_ _1046_ _1726_ VPWR VGND sg13g2_nand2_1
XFILLER_38_895 VPWR VGND sg13g2_decap_4
XFILLER_37_394 VPWR VGND sg13g2_decap_4
XFILLER_40_504 VPWR VGND sg13g2_fill_1
XFILLER_25_589 VPWR VGND sg13g2_decap_4
X_4929_ net108 VGND VPWR _0480_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\]
+ _0137_ sg13g2_dfrbpq_1
XFILLER_5_939 VPWR VGND sg13g2_decap_8
XFILLER_4_416 VPWR VGND sg13g2_decap_8
XFILLER_4_427 VPWR VGND sg13g2_fill_2
Xheichips25_bagel_21 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_0_611 VPWR VGND sg13g2_decap_8
XFILLER_48_604 VPWR VGND sg13g2_decap_8
XFILLER_47_103 VPWR VGND sg13g2_fill_2
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_48_648 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_4
XFILLER_18_61 VPWR VGND sg13g2_fill_1
XFILLER_8_722 VPWR VGND sg13g2_fill_2
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_11_261 VPWR VGND sg13g2_decap_4
XFILLER_8_799 VPWR VGND sg13g2_fill_1
XFILLER_8_788 VPWR VGND sg13g2_decap_8
XFILLER_4_950 VPWR VGND sg13g2_decap_8
X_3260_ _0994_ _0995_ _0365_ VPWR VGND sg13g2_nor2b_1
X_3191_ _0944_ _0950_ _0333_ VPWR VGND sg13g2_nor2_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_22_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_350 VPWR VGND sg13g2_fill_1
XFILLER_26_309 VPWR VGND sg13g2_decap_8
XFILLER_47_670 VPWR VGND sg13g2_fill_2
XFILLER_35_821 VPWR VGND sg13g2_fill_2
XFILLER_46_191 VPWR VGND sg13g2_decap_4
XFILLER_34_331 VPWR VGND sg13g2_decap_4
X_5058__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_34_353 VPWR VGND sg13g2_fill_2
X_2975_ _0823_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0821_ VPWR VGND
+ sg13g2_xnor2_1
X_4714_ net153 VGND VPWR _0266_ clockdiv.q2 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_30_592 VPWR VGND sg13g2_fill_1
X_4645_ net672 net723 _0198_ VPWR VGND sg13g2_nor2_1
XFILLER_30_29 VPWR VGND sg13g2_fill_2
X_4576_ net685 net736 _0129_ VPWR VGND sg13g2_nor2_1
XFILLER_2_909 VPWR VGND sg13g2_decap_8
X_3527_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\] net573 _1257_ VPWR
+ VGND sg13g2_nor2_1
X_3458_ _1173_ VPWR _1188_ VGND net547 _1187_ sg13g2_o21ai_1
X_3389_ _1119_ _1102_ _1118_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_618 VPWR VGND sg13g2_decap_8
X_5059_ net291 VGND VPWR _0606_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\]
+ _0254_ sg13g2_dfrbpq_1
XFILLER_26_898 VPWR VGND sg13g2_decap_8
XFILLER_9_519 VPWR VGND sg13g2_decap_8
XFILLER_21_581 VPWR VGND sg13g2_decap_8
XFILLER_4_202 VPWR VGND sg13g2_decap_8
XFILLER_20_62 VPWR VGND sg13g2_fill_2
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_1_986 VPWR VGND sg13g2_decap_8
X_4911__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_49_946 VPWR VGND sg13g2_decap_8
XFILLER_29_71 VPWR VGND sg13g2_decap_8
XFILLER_35_128 VPWR VGND sg13g2_fill_2
XFILLER_32_824 VPWR VGND sg13g2_decap_4
XFILLER_31_312 VPWR VGND sg13g2_decap_8
XFILLER_12_570 VPWR VGND sg13g2_decap_8
X_2760_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\] _0752_ _0482_
+ VPWR VGND sg13g2_mux2_1
X_2691_ _0738_ _0727_ _0731_ VPWR VGND sg13g2_nand2_2
X_4430_ _0643_ _1989_ _2119_ _2120_ VPWR VGND sg13g2_nor3_1
X_4361_ _2025_ _2028_ _2056_ VPWR VGND sg13g2_nor2b_1
X_4292_ _1995_ _0643_ tmds_blue.n193 VPWR VGND sg13g2_nand2_1
X_3312_ _1038_ _1014_ _1040_ _1042_ VPWR VGND sg13g2_a21o_1
X_3243_ net748 _0983_ _0984_ _0359_ VPWR VGND sg13g2_nor3_1
XFILLER_39_434 VPWR VGND sg13g2_decap_8
X_3174_ _0793_ _0939_ _0327_ VPWR VGND sg13g2_nor2_1
XFILLER_27_607 VPWR VGND sg13g2_decap_4
XFILLER_26_106 VPWR VGND sg13g2_fill_1
XFILLER_26_117 VPWR VGND sg13g2_decap_8
XFILLER_19_180 VPWR VGND sg13g2_fill_1
X_2958_ _0804_ _0792_ videogen.mem_read videogen.mem_row VPWR VGND sg13g2_a21o_2
X_2889_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\] _0782_ _0340_
+ VPWR VGND sg13g2_mux2_1
X_4628_ net688 net740 _0181_ VPWR VGND sg13g2_nor2_1
X_4559_ net682 net733 _0112_ VPWR VGND sg13g2_nor2_1
XFILLER_49_209 VPWR VGND sg13g2_decap_8
XFILLER_46_949 VPWR VGND sg13g2_decap_8
X_4865__268 VPWR VGND net268 sg13g2_tiehi
XFILLER_14_802 VPWR VGND sg13g2_fill_1
XFILLER_25_150 VPWR VGND sg13g2_fill_1
XFILLER_26_684 VPWR VGND sg13g2_fill_1
XFILLER_41_643 VPWR VGND sg13g2_fill_1
XFILLER_41_632 VPWR VGND sg13g2_decap_8
XFILLER_13_323 VPWR VGND sg13g2_fill_2
XFILLER_25_161 VPWR VGND sg13g2_decap_8
XFILLER_40_153 VPWR VGND sg13g2_fill_2
XFILLER_40_142 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_fill_2
XFILLER_14_879 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_511 VPWR VGND sg13g2_fill_1
Xoutput4 net4 tmds_clk VPWR VGND sg13g2_buf_1
XFILLER_1_783 VPWR VGND sg13g2_decap_8
XFILLER_49_765 VPWR VGND sg13g2_decap_8
XFILLER_45_971 VPWR VGND sg13g2_decap_8
X_3930_ VGND VPWR _1655_ _1656_ _1654_ _1645_ sg13g2_a21oi_2
XFILLER_17_695 VPWR VGND sg13g2_fill_1
XFILLER_32_632 VPWR VGND sg13g2_decap_8
X_3861_ VGND VPWR net616 _1584_ _1590_ _1589_ sg13g2_a21oi_1
XFILLER_20_816 VPWR VGND sg13g2_fill_1
XFILLER_32_654 VPWR VGND sg13g2_fill_2
X_3792_ _0637_ _1510_ _1521_ _1522_ VPWR VGND sg13g2_nor3_1
X_2812_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\] net764 _0765_ _0443_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_698 VPWR VGND sg13g2_fill_1
X_2743_ net762 videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\] _0748_ _0495_
+ VPWR VGND sg13g2_mux2_1
X_2674_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\] _0734_ _0559_
+ VPWR VGND sg13g2_mux2_1
X_4413_ net571 _2099_ _2103_ _0625_ VPWR VGND sg13g2_nor3_1
X_4344_ _2040_ _0844_ _2039_ VPWR VGND sg13g2_xnor2_1
X_4275_ VGND VPWR _0653_ _1954_ _1980_ _1974_ sg13g2_a21oi_1
XFILLER_39_253 VPWR VGND sg13g2_decap_8
X_3226_ VGND VPWR net610 _0970_ _0972_ videogen.fancy_shader.n646\[9\] sg13g2_a21oi_1
X_3157_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0925_ _0928_ VPWR VGND
+ sg13g2_and2_1
XFILLER_27_426 VPWR VGND sg13g2_decap_4
XFILLER_28_949 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_4
X_3088_ _0877_ _0876_ _0878_ VPWR VGND sg13g2_nor2b_2
X_4895__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_10_315 VPWR VGND sg13g2_decap_8
X_4795__384 VPWR VGND net384 sg13g2_tiehi
XFILLER_2_547 VPWR VGND sg13g2_fill_2
XFILLER_2_525 VPWR VGND sg13g2_decap_8
XFILLER_19_949 VPWR VGND sg13g2_decap_8
XFILLER_18_448 VPWR VGND sg13g2_fill_1
XFILLER_27_982 VPWR VGND sg13g2_decap_8
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_26_61 VPWR VGND sg13g2_decap_8
XFILLER_26_470 VPWR VGND sg13g2_fill_2
XFILLER_26_492 VPWR VGND sg13g2_fill_1
XFILLER_13_142 VPWR VGND sg13g2_decap_8
XFILLER_41_473 VPWR VGND sg13g2_fill_2
XFILLER_42_93 VPWR VGND sg13g2_fill_1
XFILLER_5_352 VPWR VGND sg13g2_decap_8
X_5048__157 VPWR VGND net157 sg13g2_tiehi
X_4060_ VGND VPWR _1783_ _1780_ _1769_ sg13g2_or2_1
X_3011_ net442 blue_tmds_par\[7\] net696 serialize.n429\[7\] VPWR VGND sg13g2_mux2_1
XFILLER_37_713 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_1016 VPWR VGND sg13g2_decap_8
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_36_212 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
X_4962_ net371 VGND VPWR _0509_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\]
+ _0157_ sg13g2_dfrbpq_1
XFILLER_17_470 VPWR VGND sg13g2_decap_8
X_3913_ _1639_ _1112_ _1638_ VPWR VGND sg13g2_xnor2_1
X_4893_ net210 VGND VPWR _0444_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\]
+ _0101_ sg13g2_dfrbpq_1
X_3844_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\] net566 _1573_ VPWR
+ VGND sg13g2_nor2_1
X_3775_ net597 VPWR _1505_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\]
+ net554 sg13g2_o21ai_1
X_2726_ _0707_ _0725_ _0745_ VPWR VGND sg13g2_nor2_2
X_2657_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\] _0730_ _0572_
+ VPWR VGND sg13g2_mux2_1
X_4931__100 VPWR VGND net100 sg13g2_tiehi
X_2588_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\] net772 _0700_ _0629_
+ VPWR VGND sg13g2_mux2_1
X_4327_ _2023_ net601 tmds_green.n126 VPWR VGND sg13g2_nand2_1
XFILLER_41_1000 VPWR VGND sg13g2_decap_8
X_4258_ _0883_ tmds_red.dc_balancing_reg\[2\] _0886_ _1964_ VPWR VGND sg13g2_a21o_1
X_3209_ net795 VPWR _0962_ VGND videogen.fancy_shader.n646\[2\] _0960_ sg13g2_o21ai_1
X_4189_ _1900_ _1908_ _1909_ VPWR VGND sg13g2_and2_1
XFILLER_42_226 VPWR VGND sg13g2_fill_1
XFILLER_42_204 VPWR VGND sg13g2_fill_2
XFILLER_24_974 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_fill_2
XFILLER_11_635 VPWR VGND sg13g2_fill_1
XFILLER_11_679 VPWR VGND sg13g2_fill_2
XFILLER_12_30 VPWR VGND sg13g2_decap_8
XFILLER_12_41 VPWR VGND sg13g2_fill_1
X_4717__149 VPWR VGND net149 sg13g2_tiehi
XFILLER_2_377 VPWR VGND sg13g2_decap_4
XFILLER_2_399 VPWR VGND sg13g2_decap_4
Xfanout670 net672 net670 VPWR VGND sg13g2_buf_8
XFILLER_18_201 VPWR VGND sg13g2_fill_2
Xfanout681 net682 net681 VPWR VGND sg13g2_buf_8
Xfanout692 net693 net692 VPWR VGND sg13g2_buf_8
XFILLER_46_543 VPWR VGND sg13g2_decap_4
X_5008__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_46_576 VPWR VGND sg13g2_fill_1
XFILLER_33_204 VPWR VGND sg13g2_decap_8
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_42_782 VPWR VGND sg13g2_decap_8
XFILLER_42_793 VPWR VGND sg13g2_fill_2
XFILLER_30_944 VPWR VGND sg13g2_decap_8
X_3560_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\] net556 _1290_ VPWR
+ VGND sg13g2_nor2_1
X_3491_ _1022_ _1215_ _1217_ _1218_ _1221_ VPWR VGND sg13g2_nor4_1
X_5092_ net801 VGND VPWR serialize.n428\[7\] serialize.n414\[5\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4112_ _1835_ _1833_ _1834_ VPWR VGND sg13g2_xnor2_1
X_4043_ _1761_ _1765_ _1766_ VPWR VGND sg13g2_nor2_2
X_4945_ net49 VGND VPWR _0492_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\]
+ _0149_ sg13g2_dfrbpq_1
XFILLER_24_259 VPWR VGND sg13g2_fill_1
XFILLER_21_922 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_decap_4
XFILLER_33_782 VPWR VGND sg13g2_decap_4
X_4876_ net243 VGND VPWR _0427_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\]
+ _0084_ sg13g2_dfrbpq_1
X_3827_ _1552_ _1553_ _1554_ _1555_ _1556_ VPWR VGND sg13g2_nor4_1
XFILLER_21_999 VPWR VGND sg13g2_decap_8
X_3758_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\] net574 _1488_ VPWR
+ VGND sg13g2_nor2_1
X_2709_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\] _0741_ _0531_
+ VPWR VGND sg13g2_mux2_1
X_3689_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\] net550 _1419_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_15_226 VPWR VGND sg13g2_decap_4
XFILLER_16_738 VPWR VGND sg13g2_fill_1
XFILLER_12_911 VPWR VGND sg13g2_decap_8
XFILLER_24_793 VPWR VGND sg13g2_fill_1
XFILLER_8_926 VPWR VGND sg13g2_decap_8
XFILLER_12_988 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_185 VPWR VGND sg13g2_decap_8
XFILLER_0_44 VPWR VGND sg13g2_decap_4
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_fill_2
XFILLER_0_55 VPWR VGND sg13g2_fill_1
XFILLER_19_576 VPWR VGND sg13g2_fill_1
XFILLER_0_99 VPWR VGND sg13g2_fill_1
XFILLER_22_708 VPWR VGND sg13g2_decap_8
XFILLER_34_568 VPWR VGND sg13g2_fill_1
X_2991_ VGND VPWR _0832_ _0833_ net7 _0820_ sg13g2_a21oi_1
X_4730_ net131 VGND VPWR _0281_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\]
+ _0012_ sg13g2_dfrbpq_1
XFILLER_9_64 VPWR VGND sg13g2_fill_2
X_4661_ net659 net710 _0214_ VPWR VGND sg13g2_nor2_1
X_3612_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\] net552 _1342_ VPWR
+ VGND sg13g2_nor2_1
X_4592_ net687 net738 _0145_ VPWR VGND sg13g2_nor2_1
X_3543_ _1271_ _1272_ _1273_ VPWR VGND sg13g2_nor2_1
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_3474_ VPWR _1204_ _1203_ VGND sg13g2_inv_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
XFILLER_28_29 VPWR VGND sg13g2_decap_8
X_5075_ net90 VGND VPWR _0622_ tmds_green.dc_balancing_reg\[4\] net648 sg13g2_dfrbpq_2
X_4026_ _1748_ _1735_ _1749_ VPWR VGND sg13g2_xor2_1
XFILLER_25_524 VPWR VGND sg13g2_decap_8
XFILLER_25_535 VPWR VGND sg13g2_decap_8
XFILLER_40_538 VPWR VGND sg13g2_fill_2
X_4928_ net112 VGND VPWR _0479_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\]
+ _0136_ sg13g2_dfrbpq_1
X_4859_ net280 VGND VPWR _0410_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\]
+ _0067_ sg13g2_dfrbpq_1
XFILLER_5_918 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_22 VPWR VGND uio_oe[1] sg13g2_tielo
X_4746__99 VPWR VGND net99 sg13g2_tiehi
XFILLER_0_656 VPWR VGND sg13g2_decap_8
XFILLER_28_351 VPWR VGND sg13g2_fill_2
XFILLER_11_251 VPWR VGND sg13g2_fill_2
XFILLER_11_273 VPWR VGND sg13g2_fill_2
X_5012__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_3_494 VPWR VGND sg13g2_decap_4
X_3190_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] _0948_
+ _0950_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] sg13g2_a21oi_1
XFILLER_38_115 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_fill_1
XFILLER_46_181 VPWR VGND sg13g2_decap_4
XFILLER_34_321 VPWR VGND sg13g2_decap_4
XFILLER_22_516 VPWR VGND sg13g2_fill_2
X_2974_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0821_ _0822_ VPWR VGND
+ sg13g2_and2_1
X_4713_ net154 VGND VPWR _0265_ clockdiv.q1 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
X_4644_ net664 net715 _0197_ VPWR VGND sg13g2_nor2_1
X_4575_ net676 net728 _0128_ VPWR VGND sg13g2_nor2_1
X_3526_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\] net549 _1256_ VPWR
+ VGND sg13g2_nor2_1
X_3457_ _1179_ _1186_ _1187_ VPWR VGND sg13g2_and2_1
X_3388_ _1074_ VPWR _1118_ VGND _1072_ _1075_ sg13g2_o21ai_1
X_5067__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_29_115 VPWR VGND sg13g2_fill_1
X_5058_ net306 VGND VPWR _0605_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\]
+ _0253_ sg13g2_dfrbpq_1
XFILLER_44_118 VPWR VGND sg13g2_fill_1
X_4009_ _1732_ _1084_ _1632_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_822 VPWR VGND sg13g2_fill_2
XFILLER_37_192 VPWR VGND sg13g2_decap_4
XFILLER_25_321 VPWR VGND sg13g2_fill_2
XFILLER_13_505 VPWR VGND sg13g2_decap_8
XFILLER_21_560 VPWR VGND sg13g2_decap_8
XFILLER_49_925 VPWR VGND sg13g2_decap_8
XFILLER_1_965 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_21_1020 VPWR VGND sg13g2_decap_8
XFILLER_29_94 VPWR VGND sg13g2_fill_1
XFILLER_48_479 VPWR VGND sg13g2_decap_8
XFILLER_17_822 VPWR VGND sg13g2_fill_1
XFILLER_44_641 VPWR VGND sg13g2_decap_4
XFILLER_44_630 VPWR VGND sg13g2_decap_8
XFILLER_16_332 VPWR VGND sg13g2_fill_1
XFILLER_16_354 VPWR VGND sg13g2_decap_8
XFILLER_43_184 VPWR VGND sg13g2_fill_2
XFILLER_31_335 VPWR VGND sg13g2_fill_1
XFILLER_8_531 VPWR VGND sg13g2_fill_1
X_2690_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\] _0737_ _0546_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_597 VPWR VGND sg13g2_decap_8
XFILLER_6_43 VPWR VGND sg13g2_fill_2
X_4360_ _2055_ _2041_ _2049_ VPWR VGND sg13g2_xnor2_1
X_3311_ VGND VPWR _1014_ _1038_ _1041_ _1040_ sg13g2_a21oi_1
X_4291_ VGND VPWR net606 _1993_ _0610_ _1994_ sg13g2_a21oi_1
X_3242_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\] _0814_
+ _0897_ _0984_ VPWR VGND sg13g2_and4_1
X_3173_ _0939_ net616 _0938_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_468 VPWR VGND sg13g2_decap_4
XFILLER_39_457 VPWR VGND sg13g2_fill_1
XFILLER_39_446 VPWR VGND sg13g2_decap_8
XFILLER_35_663 VPWR VGND sg13g2_fill_1
X_4949__33 VPWR VGND net33 sg13g2_tiehi
X_2957_ net429 net413 net446 serialize.n410 VPWR VGND sg13g2_nor3_2
X_2888_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\] _0782_ _0341_
+ VPWR VGND sg13g2_mux2_1
X_4627_ net688 net740 _0180_ VPWR VGND sg13g2_nor2_1
X_4558_ net689 net741 _0111_ VPWR VGND sg13g2_nor2_1
XFILLER_1_239 VPWR VGND sg13g2_fill_1
X_4489_ net653 net704 _0042_ VPWR VGND sg13g2_nor2_1
X_3509_ VGND VPWR _1235_ _1237_ _1239_ _1238_ sg13g2_a21oi_1
XFILLER_46_928 VPWR VGND sg13g2_decap_8
XFILLER_26_663 VPWR VGND sg13g2_decap_8
XFILLER_40_110 VPWR VGND sg13g2_fill_1
XFILLER_41_666 VPWR VGND sg13g2_fill_2
XFILLER_40_198 VPWR VGND sg13g2_fill_1
XFILLER_5_556 VPWR VGND sg13g2_fill_1
Xoutput5 net5 tmds_g VPWR VGND sg13g2_buf_1
XFILLER_1_762 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_fill_2
XFILLER_49_744 VPWR VGND sg13g2_decap_8
X_4844__309 VPWR VGND net309 sg13g2_tiehi
XFILLER_45_950 VPWR VGND sg13g2_decap_8
XFILLER_36_438 VPWR VGND sg13g2_fill_2
X_3860_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] VPWR _1589_ VGND net616
+ _1588_ sg13g2_o21ai_1
X_3791_ net592 _1515_ _1520_ _1521_ VPWR VGND sg13g2_nor3_1
X_2811_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\] net753 _0765_ _0444_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_165 VPWR VGND sg13g2_fill_2
X_2742_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\] _0748_ _0496_
+ VPWR VGND sg13g2_mux2_1
X_4412_ _2003_ _2100_ _2101_ _2103_ VPWR VGND sg13g2_nor3_1
XFILLER_8_394 VPWR VGND sg13g2_fill_2
X_2673_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\] _0734_ _0560_
+ VPWR VGND sg13g2_mux2_1
X_4343_ _2038_ VPWR _2039_ VGND _0847_ _2032_ sg13g2_o21ai_1
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
X_4274_ VGND VPWR _1955_ _1964_ _1979_ _1968_ sg13g2_a21oi_1
X_3225_ net747 _0971_ _0354_ VPWR VGND sg13g2_nor2_1
X_3156_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0925_ _0927_ VPWR VGND
+ sg13g2_nor2_1
XFILLER_28_928 VPWR VGND sg13g2_decap_8
X_3087_ _0870_ VPWR _0877_ VGND _0872_ _0874_ sg13g2_o21ai_1
XFILLER_42_408 VPWR VGND sg13g2_fill_1
XFILLER_36_994 VPWR VGND sg13g2_decap_8
XFILLER_23_611 VPWR VGND sg13g2_decap_8
XFILLER_22_143 VPWR VGND sg13g2_fill_2
XFILLER_35_1019 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_fill_1
X_5001__191 VPWR VGND net191 sg13g2_tiehi
X_3989_ _1714_ VPWR _1715_ VGND _1706_ _1710_ sg13g2_o21ai_1
X_4975__297 VPWR VGND net297 sg13g2_tiehi
XFILLER_19_928 VPWR VGND sg13g2_decap_8
XFILLER_46_736 VPWR VGND sg13g2_fill_1
XFILLER_45_213 VPWR VGND sg13g2_fill_2
XFILLER_26_51 VPWR VGND sg13g2_decap_4
XFILLER_27_961 VPWR VGND sg13g2_decap_8
XFILLER_14_600 VPWR VGND sg13g2_fill_1
XFILLER_14_622 VPWR VGND sg13g2_fill_2
XFILLER_42_986 VPWR VGND sg13g2_decap_8
XFILLER_41_463 VPWR VGND sg13g2_fill_2
XFILLER_14_699 VPWR VGND sg13g2_fill_1
XFILLER_42_61 VPWR VGND sg13g2_fill_1
XFILLER_9_158 VPWR VGND sg13g2_fill_2
XFILLER_42_72 VPWR VGND sg13g2_decap_8
XFILLER_6_887 VPWR VGND sg13g2_fill_1
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_fill_1
XFILLER_49_574 VPWR VGND sg13g2_decap_8
X_3010_ net418 blue_tmds_par\[6\] net695 serialize.n429\[6\] VPWR VGND sg13g2_mux2_1
XFILLER_36_268 VPWR VGND sg13g2_decap_8
XFILLER_18_994 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_4
X_4961_ net375 VGND VPWR _0508_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\]
+ _0156_ sg13g2_dfrbpq_1
X_3912_ _1638_ _1123_ _1636_ VPWR VGND sg13g2_nand2_1
X_4892_ net212 VGND VPWR _0443_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\]
+ _0100_ sg13g2_dfrbpq_1
X_3843_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\] net556 _1572_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_33_986 VPWR VGND sg13g2_decap_8
X_3774_ _1500_ _1501_ _1502_ _1503_ _1504_ VPWR VGND sg13g2_nor4_1
X_2725_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\] net790 _0744_ _0518_
+ VPWR VGND sg13g2_mux2_1
X_2656_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\] _0730_ _0573_
+ VPWR VGND sg13g2_mux2_1
X_4942__61 VPWR VGND net61 sg13g2_tiehi
X_2587_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\] net762 _0700_ _0630_
+ VPWR VGND sg13g2_mux2_1
X_4326_ net603 net601 tmds_green.n126 _2022_ VPWR VGND sg13g2_nor3_1
XFILLER_47_28 VPWR VGND sg13g2_decap_8
X_4257_ _1918_ _1959_ _1963_ VPWR VGND sg13g2_nor2_1
X_3208_ videogen.fancy_shader.n646\[2\] _0960_ _0961_ VPWR VGND sg13g2_and2_1
X_4188_ _1908_ _1907_ _1902_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_703 VPWR VGND sg13g2_fill_2
X_3139_ _0672_ VPWR _0914_ VGND videogen.mem_read _0809_ sg13g2_o21ai_1
XFILLER_28_736 VPWR VGND sg13g2_fill_1
XFILLER_28_769 VPWR VGND sg13g2_decap_4
XFILLER_24_953 VPWR VGND sg13g2_decap_8
XFILLER_35_290 VPWR VGND sg13g2_fill_1
XFILLER_11_603 VPWR VGND sg13g2_decap_4
X_5017__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_11_625 VPWR VGND sg13g2_fill_1
XFILLER_11_647 VPWR VGND sg13g2_decap_8
XFILLER_6_117 VPWR VGND sg13g2_fill_2
XFILLER_6_106 VPWR VGND sg13g2_decap_8
XFILLER_12_64 VPWR VGND sg13g2_fill_2
XFILLER_12_75 VPWR VGND sg13g2_decap_4
XFILLER_2_301 VPWR VGND sg13g2_fill_1
XFILLER_2_334 VPWR VGND sg13g2_decap_4
Xfanout660 net694 net660 VPWR VGND sg13g2_buf_8
Xfanout671 net672 net671 VPWR VGND sg13g2_buf_8
XFILLER_46_500 VPWR VGND sg13g2_decap_8
Xfanout682 net683 net682 VPWR VGND sg13g2_buf_8
Xfanout693 net694 net693 VPWR VGND sg13g2_buf_8
XFILLER_46_522 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_fill_2
XFILLER_37_50 VPWR VGND sg13g2_fill_2
XFILLER_18_235 VPWR VGND sg13g2_fill_2
XFILLER_34_717 VPWR VGND sg13g2_decap_8
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_decap_8
XFILLER_33_249 VPWR VGND sg13g2_fill_1
XFILLER_41_260 VPWR VGND sg13g2_decap_8
XFILLER_14_474 VPWR VGND sg13g2_decap_4
XFILLER_30_923 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk_regs clknet_0_clk_regs clknet_3_7__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_5015__102 VPWR VGND net102 sg13g2_tiehi
X_3490_ VPWR _1220_ _1219_ VGND sg13g2_inv_1
XFILLER_6_695 VPWR VGND sg13g2_fill_1
XFILLER_5_150 VPWR VGND sg13g2_fill_1
X_4854__290 VPWR VGND net290 sg13g2_tiehi
X_5091_ net798 VGND VPWR net428 serialize.n414\[4\] clknet_3_1__leaf_clk_regs sg13g2_dfrbpq_1
X_4111_ _1834_ _1821_ _1824_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_1018 VPWR VGND sg13g2_decap_8
X_4042_ _1762_ _1763_ _1765_ VPWR VGND sg13g2_and2_1
XFILLER_24_227 VPWR VGND sg13g2_fill_1
XFILLER_25_728 VPWR VGND sg13g2_decap_8
X_4944_ net53 VGND VPWR _0491_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\]
+ _0148_ sg13g2_dfrbpq_1
X_4875_ net245 VGND VPWR _0426_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\]
+ _0083_ sg13g2_dfrbpq_1
X_3826_ net620 VPWR _1555_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\]
+ net588 sg13g2_o21ai_1
XFILLER_20_466 VPWR VGND sg13g2_fill_2
XFILLER_21_978 VPWR VGND sg13g2_decap_8
X_3757_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\] net584 _1487_ VPWR
+ VGND sg13g2_nor2_1
X_4773__56 VPWR VGND net56 sg13g2_tiehi
X_2708_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\] _0741_ _0532_
+ VPWR VGND sg13g2_mux2_1
X_5033__279 VPWR VGND net279 sg13g2_tiehi
X_3688_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\] net573 _1418_ VPWR
+ VGND sg13g2_nor2_1
X_2639_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\] net770 _0724_ _0584_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_849 VPWR VGND sg13g2_decap_8
X_4309_ _2009_ _2001_ _2008_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_569 VPWR VGND sg13g2_fill_1
XFILLER_30_208 VPWR VGND sg13g2_decap_4
XFILLER_8_905 VPWR VGND sg13g2_decap_8
XFILLER_12_967 VPWR VGND sg13g2_decap_8
XFILLER_23_41 VPWR VGND sg13g2_fill_1
XFILLER_48_1007 VPWR VGND sg13g2_decap_8
XFILLER_3_621 VPWR VGND sg13g2_decap_8
XFILLER_2_153 VPWR VGND sg13g2_decap_4
XFILLER_19_522 VPWR VGND sg13g2_decap_8
XFILLER_19_533 VPWR VGND sg13g2_fill_2
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_46_341 VPWR VGND sg13g2_fill_1
XFILLER_19_544 VPWR VGND sg13g2_decap_8
XFILLER_0_67 VPWR VGND sg13g2_decap_4
XFILLER_19_588 VPWR VGND sg13g2_decap_8
XFILLER_0_89 VPWR VGND sg13g2_fill_1
XFILLER_34_536 VPWR VGND sg13g2_decap_4
X_2990_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\] _0829_ _0833_
+ _0819_ sg13g2_a21oi_1
XFILLER_21_219 VPWR VGND sg13g2_fill_1
XFILLER_9_43 VPWR VGND sg13g2_decap_8
X_4660_ net684 net735 _0213_ VPWR VGND sg13g2_nor2_1
XFILLER_31_1011 VPWR VGND sg13g2_decap_8
X_3611_ net593 VPWR _1341_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\]
+ net574 sg13g2_o21ai_1
X_4591_ net687 net738 _0144_ VPWR VGND sg13g2_nor2_1
X_3542_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\] net559 _1272_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_7_982 VPWR VGND sg13g2_decap_8
X_3473_ _1203_ _1201_ _1202_ VPWR VGND sg13g2_nand2_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5074_ net106 VGND VPWR _0621_ tmds_green.dc_balancing_reg\[3\] net648 sg13g2_dfrbpq_1
XFILLER_38_831 VPWR VGND sg13g2_fill_1
X_4025_ _1746_ _1747_ _1748_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_517 VPWR VGND sg13g2_decap_8
X_4927_ net116 VGND VPWR _0478_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\]
+ _0135_ sg13g2_dfrbpq_1
X_4858_ net282 VGND VPWR _0409_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\]
+ _0066_ sg13g2_dfrbpq_1
XFILLER_20_230 VPWR VGND sg13g2_fill_2
XFILLER_21_764 VPWR VGND sg13g2_fill_2
X_3809_ net598 VPWR _1539_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\]
+ net556 sg13g2_o21ai_1
X_4789_ net396 VGND VPWR _0340_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\]
+ _0040_ sg13g2_dfrbpq_1
Xheichips25_bagel_23 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_18_52 VPWR VGND sg13g2_decap_8
XFILLER_44_823 VPWR VGND sg13g2_decap_4
XFILLER_16_503 VPWR VGND sg13g2_fill_2
XFILLER_29_897 VPWR VGND sg13g2_decap_8
XFILLER_16_536 VPWR VGND sg13g2_fill_2
XFILLER_43_399 VPWR VGND sg13g2_decap_4
XFILLER_31_539 VPWR VGND sg13g2_decap_8
XFILLER_34_95 VPWR VGND sg13g2_decap_8
XFILLER_7_212 VPWR VGND sg13g2_fill_2
XFILLER_12_786 VPWR VGND sg13g2_decap_8
XFILLER_7_256 VPWR VGND sg13g2_fill_2
XFILLER_4_985 VPWR VGND sg13g2_decap_8
X_2973_ _0670_ _0683_ _0821_ VPWR VGND sg13g2_nor2_2
XFILLER_15_580 VPWR VGND sg13g2_decap_8
X_4712_ net156 VGND VPWR _0264_ tmds_blue.dc_balancing_reg\[0\] net641 sg13g2_dfrbpq_1
XFILLER_15_591 VPWR VGND sg13g2_fill_2
X_4643_ net663 net714 _0196_ VPWR VGND sg13g2_nor2_1
X_4574_ net685 net736 _0127_ VPWR VGND sg13g2_nor2_1
X_3525_ _1255_ net627 net625 VPWR VGND sg13g2_nand2b_1
X_3456_ _1184_ _1185_ _1182_ _1186_ VPWR VGND sg13g2_nand3_1
X_3387_ _1116_ _1092_ _1117_ VPWR VGND sg13g2_xor2_1
X_5057_ net345 VGND VPWR _0604_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\]
+ _0252_ sg13g2_dfrbpq_1
X_4008_ _1731_ _1076_ _1729_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_303 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_fill_1
XFILLER_5_749 VPWR VGND sg13g2_decap_8
XFILLER_0_410 VPWR VGND sg13g2_decap_8
XFILLER_1_944 VPWR VGND sg13g2_decap_8
XFILLER_20_97 VPWR VGND sg13g2_decap_8
XFILLER_49_904 VPWR VGND sg13g2_decap_8
Xhold40 serialize.n417\[5\] VPWR VGND net445 sg13g2_dlygate4sd3_1
XFILLER_16_322 VPWR VGND sg13g2_decap_4
XFILLER_45_94 VPWR VGND sg13g2_fill_1
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_12_594 VPWR VGND sg13g2_decap_8
XFILLER_6_66 VPWR VGND sg13g2_fill_2
X_3310_ _1023_ VPWR _1040_ VGND _1015_ _1024_ sg13g2_o21ai_1
X_4290_ net797 VPWR _1994_ VGND net607 hsync sg13g2_o21ai_1
XFILLER_4_793 VPWR VGND sg13g2_decap_8
X_3241_ _0983_ _0980_ videogen.fancy_shader.video_y\[3\] _0976_ videogen.fancy_shader.video_y\[2\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_39_414 VPWR VGND sg13g2_fill_2
X_3172_ _0793_ _0937_ _0938_ _0326_ VPWR VGND sg13g2_nor3_1
XFILLER_35_642 VPWR VGND sg13g2_decap_8
XFILLER_35_675 VPWR VGND sg13g2_decap_8
XFILLER_22_314 VPWR VGND sg13g2_fill_2
XFILLER_22_325 VPWR VGND sg13g2_fill_2
XFILLER_23_826 VPWR VGND sg13g2_decap_8
X_2956_ VGND VPWR _0649_ _0812_ _0003_ net747 sg13g2_a21oi_1
X_2887_ _0782_ _0702_ _0713_ VPWR VGND sg13g2_nand2_2
X_4626_ net688 net740 _0179_ VPWR VGND sg13g2_nor2_1
X_4557_ net681 net732 _0110_ VPWR VGND sg13g2_nor2_1
X_3508_ _1238_ _1232_ _1227_ VPWR VGND sg13g2_nand2b_1
X_4488_ net684 net735 _0041_ VPWR VGND sg13g2_nor2_1
X_3439_ VPWR _1169_ _1168_ VGND sg13g2_inv_1
XFILLER_46_907 VPWR VGND sg13g2_decap_8
X_5109_ net796 VGND VPWR serialize.n429\[6\] serialize.n417\[4\] clknet_3_0__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_18_609 VPWR VGND sg13g2_decap_8
XFILLER_41_623 VPWR VGND sg13g2_decap_4
XFILLER_41_601 VPWR VGND sg13g2_decap_8
XFILLER_13_325 VPWR VGND sg13g2_fill_1
XFILLER_14_826 VPWR VGND sg13g2_fill_2
XFILLER_15_31 VPWR VGND sg13g2_decap_8
XFILLER_15_42 VPWR VGND sg13g2_fill_2
XFILLER_12_1009 VPWR VGND sg13g2_decap_8
XFILLER_5_502 VPWR VGND sg13g2_decap_8
XFILLER_31_63 VPWR VGND sg13g2_fill_1
Xoutput6 net6 tmds_r VPWR VGND sg13g2_buf_1
XFILLER_1_741 VPWR VGND sg13g2_decap_8
XFILLER_49_723 VPWR VGND sg13g2_fill_2
XFILLER_0_240 VPWR VGND sg13g2_decap_4
XFILLER_0_284 VPWR VGND sg13g2_decap_8
XFILLER_0_295 VPWR VGND sg13g2_fill_2
XFILLER_29_491 VPWR VGND sg13g2_fill_2
X_5024__373 VPWR VGND net373 sg13g2_tiehi
XFILLER_44_450 VPWR VGND sg13g2_decap_8
XFILLER_16_141 VPWR VGND sg13g2_fill_1
XFILLER_17_675 VPWR VGND sg13g2_decap_8
XFILLER_32_656 VPWR VGND sg13g2_fill_1
X_5053__55 VPWR VGND net55 sg13g2_tiehi
X_3790_ _1516_ _1517_ _1518_ _1519_ _1520_ VPWR VGND sg13g2_nor4_1
X_2810_ _0721_ _0723_ _0765_ VPWR VGND sg13g2_nor2_2
XFILLER_31_144 VPWR VGND sg13g2_decap_8
XFILLER_32_689 VPWR VGND sg13g2_fill_2
X_2741_ _0748_ _0688_ _0727_ VPWR VGND sg13g2_nand2_2
XFILLER_8_373 VPWR VGND sg13g2_fill_2
XFILLER_9_896 VPWR VGND sg13g2_decap_8
X_4411_ VPWR _2102_ _2101_ VGND sg13g2_inv_1
X_2672_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\] _0734_ _0561_
+ VPWR VGND sg13g2_mux2_1
X_4342_ _2038_ _0847_ _2037_ VPWR VGND sg13g2_nand2_1
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
X_4273_ _1961_ _1977_ _1978_ VPWR VGND sg13g2_nor2_1
X_3224_ _0971_ net610 _0970_ VPWR VGND sg13g2_xnor2_1
.ends

