// A crude SRAM for testing with an initial state

module SRAM #(parameter ADR = 10, parameter DAT = 32, parameter DPTH = 1024)(
  output logic [DAT-1:0] DOUT,
  input logic [DAT-1:0] DIN,
  input logic [ADR-1:0] ADDR,
  input logic WE, RD, clk, rst_n
);

  // **************
  // Instr Mem
  // **************
  initial 
  begin
      $readmemh("image.txt", SRAMs);
  end

  //internal variables
  logic [DAT-1:0] SRAMs [DPTH-1:0];

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      SRAMs[0]   <= 32'h11111112;
      SRAMs[1]   <= 32'h22222333;
      SRAMs[2]   <= 32'h33344444;
      SRAMs[3]   <= 32'h45555555;
      SRAMs[4]   <= 32'h66666677;
      SRAMs[5]   <= 32'h77778888;
      SRAMs[6]   <= 32'h88999999;
      SRAMs[7]   <= 32'hAAAAAAAB;
      SRAMs[8]   <= 32'h11414144;
      SRAMs[9]   <= 32'h42444344;
      SRAMs[10]  <= 32'h43444444;
      SRAMs[11]  <= 32'h45444544;
      SRAMs[12]  <= 32'h46444744;
      SRAMs[13]  <= 32'h47788888;
      SRAMs[14]  <= 32'h88999999;
      SRAMs[15]  <= 32'hAAAAAABB;
      SRAMs[16]  <= 32'h14040400;
      SRAMs[17]  <= 32'h04000400;
      SRAMs[18]  <= 32'h04040400;
      SRAMs[19]  <= 32'h04000400;
      SRAMs[20]  <= 32'h04000400;
      SRAMs[21]  <= 32'h04788888;
      SRAMs[22]  <= 32'h8999999A;
      SRAMs[23]  <= 32'hAAAAAABB;
      SRAMs[24]  <= 32'h14040404;
      SRAMs[25]  <= 32'h42404404;
      SRAMs[26]  <= 32'h44040440;
      SRAMs[27]  <= 32'h44040404;
      SRAMs[28]  <= 32'h46440404;
      SRAMs[29]  <= 32'h47888888;
      SRAMs[30]  <= 32'h8999999A;
      SRAMs[31]  <= 32'hAAAAABBB;
      SRAMs[32]  <= 32'h14000400;
      SRAMs[33]  <= 32'h42404404;
      SRAMs[34]  <= 32'h34000440;
      SRAMs[35]  <= 32'h44000400;
      SRAMs[36]  <= 32'h04000400;
      SRAMs[37]  <= 32'h04888888;
      SRAMs[38]  <= 32'h999999AA;
      SRAMs[39]  <= 32'hAAAAABBB;
      SRAMs[40]  <= 32'h14040404;
      SRAMs[41]  <= 32'h42404404;
      SRAMs[42]  <= 32'h44040440;
      SRAMs[43]  <= 32'h44044644;
      SRAMs[44]  <= 32'h04044744;
      SRAMs[45]  <= 32'h04888888;
      SRAMs[46]  <= 32'h999999AA;
      SRAMs[47]  <= 32'hAAAABBBB;
      SRAMs[48]  <= 32'h14040400;
      SRAMs[49]  <= 32'h04000400;
      SRAMs[50]  <= 32'h04040400;
      SRAMs[51]  <= 32'h04045400;
      SRAMs[52]  <= 32'h04000400;
      SRAMs[53]  <= 32'h04888889;
      SRAMs[54]  <= 32'h99999AAA;
      SRAMs[55]  <= 32'hAAAABBBB;
      SRAMs[56]  <= 32'h11424244;
      SRAMs[57]  <= 32'h43444344;
      SRAMs[58]  <= 32'h44444444;
      SRAMs[59]  <= 32'h45456644;
      SRAMs[60]  <= 32'h46444744;
      SRAMs[61]  <= 32'h48888889;
      SRAMs[62]  <= 32'h99999AAA;
      SRAMs[63]  <= 32'hAAABBBBB;
      SRAMs[64]  <= 32'h11122222;
      SRAMs[65]  <= 32'h23333334;
      SRAMs[66]  <= 32'h44444555;
      SRAMs[67]  <= 32'h55556666;
      SRAMs[68]  <= 32'h66777777;
      SRAMs[69]  <= 32'h88888899;
      SRAMs[70]  <= 32'h9999AAAA;
      SRAMs[71]  <= 32'hAAABBBBB;
      SRAMs[72]  <= 32'h11222222;
      SRAMs[73]  <= 32'h33333334;
      SRAMs[74]  <= 32'h44444555;
      SRAMs[75]  <= 32'h55566666;
      SRAMs[76]  <= 32'h67777778;
      SRAMs[77]  <= 32'h88888899;
      SRAMs[78]  <= 32'h9999AAAA;
      SRAMs[79]  <= 32'hAABBBBBB;
      SRAMs[80]  <= 32'h11222222;
      SRAMs[81]  <= 32'h33333344;
      SRAMs[82]  <= 32'h44445555;
      SRAMs[83]  <= 32'h55566666;
      SRAMs[84]  <= 32'h67777778;
      SRAMs[85]  <= 32'h88888999;
      SRAMs[86]  <= 32'h999AAAAA;
      SRAMs[87]  <= 32'hAABBBBBB;
      SRAMs[88]  <= 32'h12222223;
      SRAMs[89]  <= 32'h33333344;
      SRAMs[90]  <= 32'h44445555;
      SRAMs[91]  <= 32'h55666666;
      SRAMs[92]  <= 32'h77777788;
      SRAMs[93]  <= 32'h88888999;
      SRAMs[94]  <= 32'h999AAAAA;
      SRAMs[95]  <= 32'hABBBBBBC;
      SRAMs[96]  <= 32'h12222223;
      SRAMs[97]  <= 32'h33333444;
      SRAMs[98]  <= 32'h44455555;
      SRAMs[99]  <= 32'h55666666;
      SRAMs[100] <= 32'h77777788;
      SRAMs[101] <= 32'h88889999;
      SRAMs[102] <= 32'h99AAAAAA;
      SRAMs[103] <= 32'hABBBBBBC;
      SRAMs[104] <= 32'h22222233;
      SRAMs[105] <= 32'h33333444;
      SRAMs[106] <= 32'h44455555;
      SRAMs[107] <= 32'h56666667;
      SRAMs[108] <= 32'h77777888;
      SRAMs[109] <= 32'h88889999;
      SRAMs[110] <= 32'h99AAAAAA;
      SRAMs[111] <= 32'hBBBBBBCC;
      SRAMs[112] <= 32'h22222233;
      SRAMs[113] <= 32'h33334444;
      SRAMs[114] <= 32'h44555555;
      SRAMs[115] <= 32'h56666667;
      SRAMs[116] <= 32'h77777888;
      SRAMs[117] <= 32'h88899999;
      SRAMs[118] <= 32'h9AAAAAAA;
      SRAMs[119] <= 32'hBBBBBBCC;
      SRAMs[120] <= 32'h22222333;
      SRAMs[121] <= 32'h33334444;
      SRAMs[122] <= 32'h44555555;
      SRAMs[123] <= 32'h66666677;
      SRAMs[124] <= 32'h77778888;
      SRAMs[125] <= 32'h88899999;
      SRAMs[126] <= 32'h9AAAAAAB;
      SRAMs[127] <= 32'hBBBBBCCC;
      SRAMs[128] <= 32'h22222333;
      SRAMs[129] <= 32'h33344444;
      SRAMs[130] <= 32'h45555555;
      SRAMs[131] <= 32'h66666677;
      SRAMs[132] <= 32'h77778888;
      SRAMs[133] <= 32'h88999999;
      SRAMs[134] <= 32'hAAAAAAAB;
      SRAMs[135] <= 32'hBBBBBCCC;
      SRAMs[136] <= 32'h22223333;
      SRAMs[137] <= 32'h33344444;
      SRAMs[138] <= 32'h45555556;
      SRAMs[139] <= 32'h66666777;
      SRAMs[140] <= 32'h77788888;
      SRAMs[141] <= 32'h88999999;
      SRAMs[142] <= 32'hAAAAAABB;
      SRAMs[143] <= 32'hBBBBCCCC;
      SRAMs[144] <= 32'h22223333;
      SRAMs[145] <= 32'h33444444;
      SRAMs[146] <= 32'h55555556;
      SRAMs[147] <= 32'h66666777;
      SRAMs[148] <= 32'h77788888;
      SRAMs[149] <= 32'h8999999A;
      SRAMs[150] <= 32'hAAAAAABB;
      SRAMs[151] <= 32'hBBBBCCCC;
      SRAMs[152] <= 32'h22535355;
      SRAMs[153] <= 32'h53555455;
      SRAMs[154] <= 32'h55555556;
      SRAMs[155] <= 32'h66557755;
      SRAMs[156] <= 32'h57555855;
      SRAMs[157] <= 32'h5999999A;
      SRAMs[158] <= 32'hAAAAABBB;
      SRAMs[159] <= 32'hBBBCCCCC;
      SRAMs[160] <= 32'h25050500;
      SRAMs[161] <= 32'h05000500;
      SRAMs[162] <= 32'h55000505;
      SRAMs[163] <= 32'h65005500;
      SRAMs[164] <= 32'h05000500;
      SRAMs[165] <= 32'h059999AA;
      SRAMs[166] <= 32'hAAAAABBB;
      SRAMs[167] <= 32'hBBBCCCCC;
      SRAMs[168] <= 32'h25050505;
      SRAMs[169] <= 32'h54505505;
      SRAMs[170] <= 32'h05055505;
      SRAMs[171] <= 32'h65050505;
      SRAMs[172] <= 32'h55050505;
      SRAMs[173] <= 32'h599999AA;
      SRAMs[174] <= 32'hAAAABBBB;
      SRAMs[175] <= 32'hBBCCCCCC;
      SRAMs[176] <= 32'h25000500;
      SRAMs[177] <= 32'h54505505;
      SRAMs[178] <= 32'h05005505;
      SRAMs[179] <= 32'h65005500;
      SRAMs[180] <= 32'h55000505;
      SRAMs[181] <= 32'h05999AAA;
      SRAMs[182] <= 32'hAAAABBBB;
      SRAMs[183] <= 32'hBBCCCCCC;
      SRAMs[184] <= 32'h25050505;
      SRAMs[185] <= 32'h54505505;
      SRAMs[186] <= 32'h05055505;
      SRAMs[187] <= 32'h55050505;
      SRAMs[188] <= 32'h55005505;
      SRAMs[189] <= 32'h05999AAA;
      SRAMs[190] <= 32'hAAABBBBB;
      SRAMs[191] <= 32'hBCCCCCCC;
      SRAMs[192] <= 32'h25050500;
      SRAMs[193] <= 32'h05000500;
      SRAMs[194] <= 32'h55000500;
      SRAMs[195] <= 32'h05005500;
      SRAMs[196] <= 32'h05050500;
      SRAMs[197] <= 32'h0599AAAA;
      SRAMs[198] <= 32'hAAABBBBB;
      SRAMs[199] <= 32'hBCCCCCCD;
      SRAMs[200] <= 32'h33535355;
      SRAMs[201] <= 32'h54555555;
      SRAMs[202] <= 32'h55555655;
      SRAMs[203] <= 32'h57557755;
      SRAMs[204] <= 32'h58585855;
      SRAMs[205] <= 32'h5999AAAA;
      SRAMs[206] <= 32'hAABBBBBB;
      SRAMs[207] <= 32'hCCCCCCCD;
      SRAMs[208] <= 32'h33333344;
      SRAMs[209] <= 32'h44445555;
      SRAMs[210] <= 32'h55566666;
      SRAMs[211] <= 32'h67777778;
      SRAMs[212] <= 32'h88888999;
      SRAMs[213] <= 32'h999AAAAA;
      SRAMs[214] <= 32'hAABBBBBB;
      SRAMs[215] <= 32'hCCCCCCDD;
      SRAMs[216] <= 32'h33333344;
      SRAMs[217] <= 32'h44445555;
      SRAMs[218] <= 32'h55666666;
      SRAMs[219] <= 32'h77777788;
      SRAMs[220] <= 32'h88888999;
      SRAMs[221] <= 32'h999AAAAA;
      SRAMs[222] <= 32'hABBBBBBC;
      SRAMs[223] <= 32'hCCCCCCDD;
      SRAMs[224] <= 32'h33333444;
      SRAMs[225] <= 32'h44455555;
      SRAMs[226] <= 32'h55666666;
      SRAMs[227] <= 32'h77777788;
      SRAMs[228] <= 32'h88889999;
      SRAMs[229] <= 32'h99AAAAAA;
      SRAMs[230] <= 32'hABBBBBBC;
      SRAMs[231] <= 32'hCCCCCDDD;
      SRAMs[232] <= 32'h33333444;
      SRAMs[233] <= 32'h44455555;
      SRAMs[234] <= 32'h56666667;
      SRAMs[235] <= 32'h77777888;
      SRAMs[236] <= 32'h88889999;
      SRAMs[237] <= 32'h99AAAAAA;
      SRAMs[238] <= 32'hBBBBBBCC;
      SRAMs[239] <= 32'hCCCCCDDD;
      SRAMs[240] <= 32'h33334444;
      SRAMs[241] <= 32'h44555555;
      SRAMs[242] <= 32'h56666667;
      SRAMs[243] <= 32'h77777888;
      SRAMs[244] <= 32'h88899999;
      SRAMs[245] <= 32'h9AAAAAAA;
      SRAMs[246] <= 32'hBBBBBBCC;
      SRAMs[247] <= 32'hCCCCDDDD;
      SRAMs[248] <= 32'h33334444;
      SRAMs[249] <= 32'h44555555;
      SRAMs[250] <= 32'h66666677;
      SRAMs[251] <= 32'h77778888;
      SRAMs[252] <= 32'h88899999;
      SRAMs[253] <= 32'h9AAAAAAB;
      SRAMs[254] <= 32'hBBBBBCCC;
      SRAMs[255] <= 32'hCCCCDDDD;
      SRAMs[256] <= 32'h33344444;
      SRAMs[257] <= 32'h45555555;
      SRAMs[258] <= 32'h66666677;
      SRAMs[259] <= 32'h77778888;
      SRAMs[260] <= 32'h88999999;
      SRAMs[261] <= 32'hAAAAAAAB;
      SRAMs[262] <= 32'hBBBBBCCC;
      SRAMs[263] <= 32'hCCCDDDDD;
      SRAMs[264] <= 32'h33222444;
      SRAMs[265] <= 32'h45222556;
      SRAMs[266] <= 32'h66222727;
      SRAMs[267] <= 32'h27222888;
      SRAMs[268] <= 32'h88222922;
      SRAMs[269] <= 32'h2AAAAABB;
      SRAMs[270] <= 32'hBBBBCCCC;
      SRAMs[271] <= 32'hCCCDDDDD;
      SRAMs[272] <= 32'h32000244;
      SRAMs[273] <= 32'h52000256;
      SRAMs[274] <= 32'h62000202;
      SRAMs[275] <= 32'h02000288;
      SRAMs[276] <= 32'h82000200;
      SRAMs[277] <= 32'h02AAAABB;
      SRAMs[278] <= 32'hBBBBCCCC;
      SRAMs[279] <= 32'hCCDDDDDD;
      SRAMs[280] <= 32'h33220222;
      SRAMs[281] <= 32'h22020266;
      SRAMs[282] <= 32'h62020202;
      SRAMs[283] <= 32'h02022888;
      SRAMs[284] <= 32'h89220202;
      SRAMs[285] <= 32'h2AAAABBB;
      SRAMs[286] <= 32'hBBBCCCCC;
      SRAMs[287] <= 32'hCCDDDDDD;
      SRAMs[288] <= 32'h32000200;
      SRAMs[289] <= 32'h02000266;
      SRAMs[290] <= 32'h62000202;
      SRAMs[291] <= 32'h02020288;
      SRAMs[292] <= 32'h92000200;
      SRAMs[293] <= 32'h02AAABBB;
      SRAMs[294] <= 32'hBBBCCCCC;
      SRAMs[295] <= 32'hCDDDDDDE;
      SRAMs[296] <= 32'h34220222;
      SRAMs[297] <= 32'h22020266;
      SRAMs[298] <= 32'h62020202;
      SRAMs[299] <= 32'h02020288;
      SRAMs[300] <= 32'h92022922;
      SRAMs[301] <= 32'h02AABBBB;
      SRAMs[302] <= 32'hBBCCCCCC;
      SRAMs[303] <= 32'hCDDDDDDE;
      SRAMs[304] <= 32'h42000255;
      SRAMs[305] <= 32'h52000266;
      SRAMs[306] <= 32'h62020200;
      SRAMs[307] <= 32'h02000289;
      SRAMs[308] <= 32'h92000200;
      SRAMs[309] <= 32'h02AABBBB;
      SRAMs[310] <= 32'hBBCCCCCC;
      SRAMs[311] <= 32'hDDDDDDEE;
      SRAMs[312] <= 32'h44222455;
      SRAMs[313] <= 32'h55222666;
      SRAMs[314] <= 32'h66272722;
      SRAMs[315] <= 32'h28222889;
      SRAMs[316] <= 32'h99222A22;
      SRAMs[317] <= 32'h2AABBBBB;
      SRAMs[318] <= 32'hBCCCCCCC;
      SRAMs[319] <= 32'hDDDDDDEE;
      SRAMs[320] <= 32'h44444555;
      SRAMs[321] <= 32'h55556666;
      SRAMs[322] <= 32'h66777777;
      SRAMs[323] <= 32'h88888899;
      SRAMs[324] <= 32'h9999AAAA;
      SRAMs[325] <= 32'hAAABBBBB;
      SRAMs[326] <= 32'hBCCCCCCD;
      SRAMs[327] <= 32'hDDDDDEEE;
      SRAMs[328] <= 32'h44444555;
      SRAMs[329] <= 32'h55566666;
      SRAMs[330] <= 32'h67777778;
      SRAMs[331] <= 32'h88888899;
      SRAMs[332] <= 32'h9999AAAA;
      SRAMs[333] <= 32'hAABBBBBB;
      SRAMs[334] <= 32'hCCCCCCCD;
      SRAMs[335] <= 32'hDDDDDEEE;
      SRAMs[336] <= 32'h44445555;
      SRAMs[337] <= 32'h55566666;
      SRAMs[338] <= 32'h67777778;
      SRAMs[339] <= 32'h88888999;
      SRAMs[340] <= 32'h999AAAAA;
      SRAMs[341] <= 32'hAABBBBBB;
      SRAMs[342] <= 32'hCCCCCCDD;
      SRAMs[343] <= 32'hDDDDEEEE;
      SRAMs[344] <= 32'h44445555;
      SRAMs[345] <= 32'h55666666;
      SRAMs[346] <= 32'h77777788;
      SRAMs[347] <= 32'h88888999;
      SRAMs[348] <= 32'h999AAAAA;
      SRAMs[349] <= 32'hABBBBBBC;
      SRAMs[350] <= 32'hCCCCCCDD;
      SRAMs[351] <= 32'hDDDDEEEE;
      SRAMs[352] <= 32'h44455555;
      SRAMs[353] <= 32'h55666666;
      SRAMs[354] <= 32'h77777788;
      SRAMs[355] <= 32'h88889999;
      SRAMs[356] <= 32'h99AAAAAA;
      SRAMs[357] <= 32'hABBBBBBC;
      SRAMs[358] <= 32'hCCCCCDDD;
      SRAMs[359] <= 32'hDDDEEEEE;
      SRAMs[360] <= 32'h44455555;
      SRAMs[361] <= 32'h56666667;
      SRAMs[362] <= 32'h77777888;
      SRAMs[363] <= 32'h88889999;
      SRAMs[364] <= 32'h99AAAAAA;
      SRAMs[365] <= 32'hBBBBBBCC;
      SRAMs[366] <= 32'hCCCCCDDD;
      SRAMs[367] <= 32'hDDDEEEEE;
      SRAMs[368] <= 32'h44555555;
      SRAMs[369] <= 32'h56666667;
      SRAMs[370] <= 32'h77777888;
      SRAMs[371] <= 32'h88899999;
      SRAMs[372] <= 32'h9AAAAAAA;
      SRAMs[373] <= 32'hBBBBBBCC;
      SRAMs[374] <= 32'hCCCCDDDD;
      SRAMs[375] <= 32'hDDEEEEEE;
      SRAMs[376] <= 32'h44555555;
      SRAMs[377] <= 32'h66666677;
      SRAMs[378] <= 32'h77778888;
      SRAMs[379] <= 32'h88899999;
      SRAMs[380] <= 32'h9AAAAAAB;
      SRAMs[381] <= 32'hBBBBBCCC;
      SRAMs[382] <= 32'hCCCCDDDD;
      SRAMs[383] <= 32'hDDEEEEEE;
      
      //SRAMs[0:383] <= {32'h11111112, 32'h22222333, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'h11414144, 32'h42444344, 32'h43444444, 32'h45444544, 32'h46444777, 32'h77788888, 32'h88999999, 32'hAAAAAABB, 32'h14040400, 32'h04000400, 32'h04040400, 32'h04000400, 32'h04000477, 32'h77788888, 32'h8999999A, 32'hAAAAAABB, 32'h14040404, 32'h42404404, 32'h44040440, 32'h44040404, 32'h46440477, 32'h77888888, 32'h8999999A, 32'hAAAAABBB, 32'h14000400, 32'h42404404, 32'h34000440, 32'h44000400, 32'h04000477, 32'h77888888, 32'h999999AA, 32'hAAAAABBB, 32'h14040404, 32'h42404404, 32'h44040440, 32'h44044644, 32'h04044777, 32'h78888888, 32'h999999AA, 32'hAAAABBBB, 32'h14040400, 32'h04000400, 32'h04040400, 32'h04045400, 32'h04000477, 32'h78888889, 32'h99999AAA, 32'hAAAABBBB, 32'h11424244, 32'h43444344, 32'h44444444, 32'h45456644, 32'h46444777, 32'h88888889, 32'h99999AAA, 32'hAAABBBBB, 32'h11122222, 32'h23333334, 32'h44444555, 32'h55556666, 32'h66777777, 32'h88888899, 32'h9999AAAA, 32'hAAABBBBB, 32'h11222222, 32'h33333334, 32'h44444555, 32'h55566666, 32'h67777778, 32'h88888899, 32'h9999AAAA, 32'hAABBBBBB, 32'h11222222, 32'h33333344, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'h12222223, 32'h33333344, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'h12222223, 32'h33333444, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'h22222233, 32'h33333444, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'h22222233, 32'h33334444, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'h22222333, 32'h33334444, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'h22222333, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'hBBBBBCCC, 32'h22223333, 32'h33344444, 32'h45555556, 32'h66666777, 32'h77788888, 32'h88999999, 32'hAAAAAABB, 32'hBBBBCCCC, 32'h22223333, 32'h33444444, 32'h55555556, 32'h66666777, 32'h77788888, 32'h8999999A, 32'hAAAAAABB, 32'hBBBBCCCC, 32'h22535355, 32'h53555455, 32'h55555556, 32'h66557755, 32'h57555855, 32'h5999999A, 32'hAAAAABBB, 32'hBBBCCCCC, 32'h25050500, 32'h05000500, 32'h55000505, 32'h65005500, 32'h05000500, 32'h059999AA, 32'hAAAAABBB, 32'hBBBCCCCC, 32'h25050505, 32'h54505505, 32'h05055505, 32'h65050505, 32'h55050505, 32'h599999AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'h25000500, 32'h54505505, 32'h05005505, 32'h65005500, 32'h55000505, 32'h05999AAA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'h25050505, 32'h54505505, 32'h05055505, 32'h55050505, 32'h55005505, 32'h05999AAA, 32'hAAABBBBB, 32'hBCCCCCCC, 32'h25050500, 32'h05000500, 32'h55000500, 32'h05005500, 32'h05050500, 32'h0599AAAA, 32'hAAABBBBB, 32'hBCCCCCCD, 32'h33535355, 32'h54555555, 32'h55555655, 32'h57557755, 32'h58585855, 32'h5999AAAA, 32'hAABBBBBB, 32'hCCCCCCCD, 32'h33333344, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'hCCCCCCDD, 32'h33333344, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'hCCCCCCDD, 32'h33333444, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'hCCCCCDDD, 32'h33333444, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'hCCCCCDDD, 32'h33334444, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'hCCCCDDDD, 32'h33334444, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'hCCCCDDDD, 32'h33344444, 32'h45555555, 32'h66666677, 32'h77778888, 32'h88999999, 32'hAAAAAAAB, 32'hBBBBBCCC, 32'hCCCDDDDD, 32'h33222444, 32'h45222556, 32'h66222727, 32'h27222888, 32'h88222999, 32'hAAAAAABB, 32'hBBBBCCCC, 32'hCCCDDDDD, 32'h32000244, 32'h52000256, 32'h62000202, 32'h02000288, 32'h8200029A, 32'hAAAAAABB, 32'hBBBBCCCC, 32'hCCDDDDDD, 32'h33220222, 32'h22020266, 32'h62020202, 32'h02022888, 32'h8922029A, 32'hAAAAABBB, 32'hBBBCCCCC, 32'hCCDDDDDD, 32'h32000200, 32'h02000266, 32'h62000202, 32'h02020288, 32'h920002AA, 32'hAAAAABBB, 32'hBBBCCCCC, 32'hCDDDDDDE, 32'h34220222, 32'h22020266, 32'h62020202, 32'h02020288, 32'h920229AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'hCDDDDDDE, 32'h42000255, 32'h52000266, 32'h62020200, 32'h02000289, 32'h920002AA, 32'hAAAABBBB, 32'hBBCCCCCC, 32'hDDDDDDEE, 32'h44222455, 32'h55222666, 32'h66272722, 32'h28222889, 32'h99222AAA, 32'hAAABBBBB, 32'hBCCCCCCC, 32'hDDDDDDEE, 32'h44444555, 32'h55556666, 32'h66777777, 32'h88888899, 32'h9999AAAA, 32'hAAABBBBB, 32'hBCCCCCCD, 32'hDDDDDEEE, 32'h44444555, 32'h55566666, 32'h67777778, 32'h88888899, 32'h9999AAAA, 32'hAABBBBBB, 32'hCCCCCCCD, 32'hDDDDDEEE, 32'h44445555, 32'h55566666, 32'h67777778, 32'h88888999, 32'h999AAAAA, 32'hAABBBBBB, 32'hCCCCCCDD, 32'hDDDDEEEE, 32'h44445555, 32'h55666666, 32'h77777788, 32'h88888999, 32'h999AAAAA, 32'hABBBBBBC, 32'hCCCCCCDD, 32'hDDDDEEEE, 32'h44455555, 32'h55666666, 32'h77777788, 32'h88889999, 32'h99AAAAAA, 32'hABBBBBBC, 32'hCCCCCDDD, 32'hDDDEEEEE, 32'h44455555, 32'h56666667, 32'h77777888, 32'h88889999, 32'h99AAAAAA, 32'hBBBBBBCC, 32'hCCCCCDDD, 32'hDDDEEEEE, 32'h44555555, 32'h56666667, 32'h77777888, 32'h88899999, 32'h9AAAAAAA, 32'hBBBBBBCC, 32'hCCCCDDDD, 32'hDDEEEEEE, 32'h44555555, 32'h66666677, 32'h77778888, 32'h88899999, 32'h9AAAAAAB, 32'hBBBBBCCC, 32'hCCCCDDDD, 32'hDDEEEEEE};
    end
    else if (WE == 1'b1 && RD == 1'b0) SRAMs[ADDR] <= DIN;
    else;
  end

  assign DOUT = SRAMs[ADDR];

endmodule



