module pixel_feeder(
  input logic clk_25, rst_n,

  output logic [3:0] pixel_out,
  input logic [3:0] pixel_in,

  // Address pins
  output logic bank,
  output logic [8:0] addr,
  output logic [2:0] pix_sel,
  
  input logic disp_active, line_end, frame_end
);
  assign bank = 0;                    // Pin bank to 0 for the moment

  logic [3:0] row [5:0];              // 64-pixel buffer to hold an entire row
  logic [3:0] h_counter, v_counter;   // Counters for tracking the /10 for H and V.
  logic [5:0] h_pix, v_pix;           // Local pixel counts
  
  
  always_comb begin
    pixel_out = row[h_pix];            // Grab the specific pixel for the row
  end
  
  // Pixel Fetcher state machine
  // If we are at v_counter 9, we want to read the pixel for the next row into the buffer when h_counter gets to 9
  // We can get away with one state for reading memory as memory is running at 126 MHz while this is running at 25 MHz,
  // So memory will be ready on the negative clock edge...
  enum {idle = 0, mem_read} state, next_state;
  
  always_comb begin
    if (state == mem_read) begin
      if (h_pix == 0) {addr,pix_sel} = {(v_pix),63};                // We end up reading the last pixel of the current line at the start of the line
      else if (v_pix == 48) {addr,pix_sel} = {6'b000000,h_pix}-1;   // Edge case if we are on the last line
      else {addr,pix_sel} = {(v_pix+1),h_pix}-1;      // Set the memory address to get the nextrow
      
      next_state = idle;
    end
    else begin
      if((v_counter == 9) && (h_counter == 9) && disp_active) next_state = mem_read;
      //{addr,pix_sel} = '0;              // Clear the memory address
    end
  end

  always_ff @(posedge clk_25) begin
    if(!rst_n) state <= idle;
    else state <= next_state;
  end

  always_ff @(negedge clk_25) begin
    if(state == mem_read) begin
      // Save the pixel from the memory interface.
      if(h_pix == 0) row[63] <= pixel_in;
      else row[h_pix-1] <= pixel_in;
    end
  end
  

  // The counters that make it all work:  
  // Horizontal pixel counter. Increments every 10th pixel
  always_ff @(posedge clk_25) begin
    if (!disp_active || !rst_n) begin 
        h_counter <= 9;                // Hold at 9 during display inactive to resync.
        h_pix <= 63;                    // Hold horizontal pixel count at 63 during display inactive to resync.
    end
    if (disp_active) begin              // Only increment if the display is active
      if (h_counter < 9) h_counter <= h_counter + 1;
      else begin
        h_counter <= 0;                 
        h_pix <= h_pix + 1;             // Increment the horizontal pixel co-ordinate.
      end
    end
  end
  
  // Vertical pixel count, incremented on line_end. Async reset on frame_end
  always_ff @(posedge line_end or posedge frame_end) begin   
    if (frame_end || !rst_n) begin
      v_counter <= 9;     // resync counter on frame end
      v_pix <= 0;
    end
    else if (v_counter < 9) v_counter <= v_counter + 1;
    else begin 
      v_counter <= 0;
      if (v_pix < 47) v_pix <= v_pix +1;              // Increment the vertical pixel co-ordinate
      else v_pix <= 0;
    end
  end    
  
endmodule