* NGSPICE file created from heichips25_bagel.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

.subckt heichips25_bagel VGND VPWR clk ena rst_n tmds_b tmds_clk tmds_g tmds_r ui_in[0]
+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1]
+ uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_277 VPWR VGND sg13g2_decap_8
X_3155_ VPWR _0884_ _0883_ VGND sg13g2_inv_1
XFILLER_28_929 VPWR VGND sg13g2_decap_8
X_3086_ net427 blue_tmds_par\[5\] net694 serialize.n429\[5\] VPWR VGND sg13g2_mux2_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
XFILLER_23_623 VPWR VGND sg13g2_decap_4
XFILLER_22_133 VPWR VGND sg13g2_decap_8
XFILLER_35_494 VPWR VGND sg13g2_decap_4
X_3988_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\] net564 _1656_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_10_317 VPWR VGND sg13g2_decap_4
X_2939_ net764 _0786_ _0787_ VPWR VGND sg13g2_nor2_1
X_4609_ net655 net702 _0039_ VPWR VGND sg13g2_nor2_1
XFILLER_7_7 VPWR VGND sg13g2_fill_1
XFILLER_27_984 VPWR VGND sg13g2_decap_8
XFILLER_14_645 VPWR VGND sg13g2_fill_1
XFILLER_42_987 VPWR VGND sg13g2_decap_8
XFILLER_41_475 VPWR VGND sg13g2_fill_1
XFILLER_41_464 VPWR VGND sg13g2_fill_1
Xclkbuf_3_6__f_clk_regs clknet_0_clk_regs clknet_3_6__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_42_40 VPWR VGND sg13g2_fill_1
XFILLER_41_486 VPWR VGND sg13g2_decap_4
XFILLER_13_177 VPWR VGND sg13g2_decap_4
XFILLER_10_895 VPWR VGND sg13g2_decap_8
XFILLER_5_365 VPWR VGND sg13g2_decap_8
XFILLER_1_571 VPWR VGND sg13g2_fill_2
X_5048__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
XFILLER_49_597 VPWR VGND sg13g2_decap_8
XFILLER_37_726 VPWR VGND sg13g2_decap_4
XFILLER_36_203 VPWR VGND sg13g2_fill_1
XFILLER_18_940 VPWR VGND sg13g2_decap_8
XFILLER_36_247 VPWR VGND sg13g2_fill_1
XFILLER_33_910 VPWR VGND sg13g2_decap_8
X_4960_ net324 VGND VPWR _0388_ red_tmds_par\[9\] net641 sg13g2_dfrbpq_1
X_4891_ net68 VGND VPWR _0319_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\]
+ net631 sg13g2_dfrbpq_1
X_3911_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\] net568 _1580_ VPWR
+ VGND sg13g2_nor2_1
X_3842_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\] net565 _1511_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_453 VPWR VGND sg13g2_fill_1
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_32_486 VPWR VGND sg13g2_decap_8
XFILLER_32_497 VPWR VGND sg13g2_fill_2
XFILLER_34_1020 VPWR VGND sg13g2_decap_8
X_3773_ _1441_ VPWR _1442_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\]
+ net553 sg13g2_o21ai_1
X_2724_ _0733_ net546 _0718_ VPWR VGND sg13g2_nand2_2
X_2655_ _0700_ _0707_ _0708_ VPWR VGND sg13g2_nor2_2
X_2586_ _0642_ videogen.fancy_shader.n646\[7\] VPWR VGND sg13g2_inv_2
X_4325_ VGND VPWR net606 _1981_ _0384_ net747 sg13g2_a21oi_1
X_4256_ _1918_ _1917_ _1905_ VPWR VGND sg13g2_nand2b_1
X_3207_ _0814_ _0927_ _0303_ VPWR VGND sg13g2_nor2_1
X_4187_ _1848_ _1845_ _1840_ _1849_ VPWR VGND sg13g2_a21o_2
X_3138_ _0867_ tmds_red.n114 tmds_red.n132 VPWR VGND sg13g2_nand2_1
X_3069_ serialize.n461 serialize.n459 clknet_1_0__leaf_clk net4 VPWR VGND sg13g2_mux2_1
XFILLER_35_291 VPWR VGND sg13g2_fill_2
XFILLER_24_976 VPWR VGND sg13g2_decap_8
XFILLER_7_619 VPWR VGND sg13g2_fill_1
XFILLER_3_836 VPWR VGND sg13g2_decap_8
XFILLER_2_302 VPWR VGND sg13g2_decap_8
Xfanout650 net651 net650 VPWR VGND sg13g2_buf_8
Xfanout694 net695 net694 VPWR VGND sg13g2_buf_8
XFILLER_19_704 VPWR VGND sg13g2_decap_8
XFILLER_19_715 VPWR VGND sg13g2_fill_1
Xfanout672 net693 net672 VPWR VGND sg13g2_buf_8
Xfanout661 net662 net661 VPWR VGND sg13g2_buf_1
Xfanout683 net687 net683 VPWR VGND sg13g2_buf_8
XFILLER_46_512 VPWR VGND sg13g2_decap_8
XFILLER_18_225 VPWR VGND sg13g2_decap_4
XFILLER_46_556 VPWR VGND sg13g2_decap_8
XFILLER_19_759 VPWR VGND sg13g2_fill_2
XFILLER_15_954 VPWR VGND sg13g2_decap_8
XFILLER_42_751 VPWR VGND sg13g2_decap_8
XFILLER_41_250 VPWR VGND sg13g2_decap_8
XFILLER_30_924 VPWR VGND sg13g2_decap_8
XFILLER_5_173 VPWR VGND sg13g2_fill_2
X_5090_ net353 VGND VPWR _0514_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\]
+ _0162_ sg13g2_dfrbpq_1
XFILLER_2_880 VPWR VGND sg13g2_decap_8
X_4110_ _1759_ _1774_ _1775_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
X_4041_ _1706_ _0995_ _1192_ VPWR VGND sg13g2_nand2_2
XFILLER_49_383 VPWR VGND sg13g2_decap_8
XFILLER_25_707 VPWR VGND sg13g2_decap_8
XFILLER_18_792 VPWR VGND sg13g2_decap_8
X_4943_ net341 VGND VPWR _0371_ display_enable net636 sg13g2_dfrbpq_1
X_4874_ net94 VGND VPWR _0302_ videogen.fancy_shader.video_x\[3\] net632 sg13g2_dfrbpq_2
XFILLER_21_957 VPWR VGND sg13g2_decap_8
X_3825_ _1447_ _1493_ net2 _1494_ VPWR VGND sg13g2_nand3_1
X_3756_ _1425_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
X_2707_ _0647_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] net619 _0728_
+ VPWR VGND _0704_ sg13g2_nand4_1
X_3687_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\] net568 _1356_ VPWR
+ VGND sg13g2_nor2_1
X_2638_ _0691_ _0685_ _0690_ VPWR VGND sg13g2_nand2_2
XFILLER_0_817 VPWR VGND sg13g2_decap_8
X_4308_ _0662_ _1967_ _1968_ _1969_ _1970_ VPWR VGND sg13g2_or4_1
XFILLER_47_309 VPWR VGND sg13g2_fill_1
X_4239_ _1901_ _1073_ _1870_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_718 VPWR VGND sg13g2_fill_1
XFILLER_43_548 VPWR VGND sg13g2_decap_8
XFILLER_24_751 VPWR VGND sg13g2_fill_1
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_23_31 VPWR VGND sg13g2_fill_1
XFILLER_11_467 VPWR VGND sg13g2_decap_4
XFILLER_20_990 VPWR VGND sg13g2_decap_8
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_644 VPWR VGND sg13g2_fill_2
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_fill_2
XFILLER_0_79 VPWR VGND sg13g2_decap_4
XFILLER_34_548 VPWR VGND sg13g2_fill_1
XFILLER_21_209 VPWR VGND sg13g2_decap_4
XFILLER_30_765 VPWR VGND sg13g2_fill_1
X_4590_ net686 net738 _0020_ VPWR VGND sg13g2_nor2_1
X_3610_ _1276_ _1268_ _1278_ _1279_ VPWR VGND sg13g2_a21o_1
XFILLER_31_1012 VPWR VGND sg13g2_decap_8
X_3541_ _1187_ _1178_ _1210_ VPWR VGND sg13g2_xor2_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
X_3472_ _1116_ _1117_ _1120_ _1141_ VPWR VGND sg13g2_or3_1
X_5211_ net803 VGND VPWR serialize.n428\[3\] serialize.n414\[1\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_43_2 VPWR VGND sg13g2_fill_1
X_5142_ net61 VGND VPWR _0566_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\]
+ _0214_ sg13g2_dfrbpq_1
X_5073_ net31 VGND VPWR _0497_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\]
+ _0154_ sg13g2_dfrbpq_1
X_4024_ VGND VPWR _1667_ _1691_ _1692_ _0661_ sg13g2_a21oi_1
XFILLER_25_504 VPWR VGND sg13g2_decap_8
XFILLER_25_559 VPWR VGND sg13g2_decap_8
XFILLER_40_518 VPWR VGND sg13g2_decap_8
X_4926_ net370 VGND VPWR _0354_ videogen.fancy_shader.n646\[8\] net632 sg13g2_dfrbpq_1
X_4857_ net125 VGND VPWR _0285_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\]
+ _0016_ sg13g2_dfrbpq_1
XFILLER_21_776 VPWR VGND sg13g2_fill_1
X_3808_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\] net578 _1477_ VPWR
+ VGND sg13g2_nor2_1
X_4788_ net690 net742 _0218_ VPWR VGND sg13g2_nor2_1
XFILLER_5_909 VPWR VGND sg13g2_decap_8
XFILLER_20_286 VPWR VGND sg13g2_fill_1
XFILLER_20_297 VPWR VGND sg13g2_decap_8
X_3739_ _1407_ VPWR _1408_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\]
+ net581 sg13g2_o21ai_1
Xheichips25_bagel_24 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_28_320 VPWR VGND sg13g2_decap_4
XFILLER_29_865 VPWR VGND sg13g2_fill_1
XFILLER_18_64 VPWR VGND sg13g2_fill_1
XFILLER_29_887 VPWR VGND sg13g2_fill_2
XFILLER_43_367 VPWR VGND sg13g2_fill_1
XFILLER_43_389 VPWR VGND sg13g2_fill_1
XFILLER_8_725 VPWR VGND sg13g2_fill_2
XFILLER_8_714 VPWR VGND sg13g2_decap_8
XFILLER_4_953 VPWR VGND sg13g2_decap_8
XFILLER_3_463 VPWR VGND sg13g2_fill_1
XFILLER_3_496 VPWR VGND sg13g2_fill_1
XFILLER_39_618 VPWR VGND sg13g2_fill_2
XFILLER_46_194 VPWR VGND sg13g2_decap_8
XFILLER_46_172 VPWR VGND sg13g2_fill_2
XFILLER_34_345 VPWR VGND sg13g2_decap_4
X_2972_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\] _0795_ _0311_
+ VPWR VGND sg13g2_mux2_1
XFILLER_34_378 VPWR VGND sg13g2_fill_2
X_4711_ net681 net730 _0141_ VPWR VGND sg13g2_nor2_1
X_4642_ net665 net717 _0072_ VPWR VGND sg13g2_nor2_1
XFILLER_30_573 VPWR VGND sg13g2_decap_8
X_4573_ _2183_ _2200_ _2201_ VPWR VGND sg13g2_nor2_1
X_3524_ _1193_ _1192_ _1016_ VPWR VGND sg13g2_nand2b_1
X_3455_ VGND VPWR videogen.fancy_shader.n646\[7\] net629 _1124_ _1123_ sg13g2_a21oi_1
X_3386_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[3\] _1055_ _0369_ _1056_
+ sg13g2_a21oi_1
X_5125_ net189 VGND VPWR _0549_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\]
+ _0197_ sg13g2_dfrbpq_1
XFILLER_38_640 VPWR VGND sg13g2_decap_8
X_5056_ net84 VGND VPWR _0484_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\]
+ _0141_ sg13g2_dfrbpq_1
XFILLER_29_139 VPWR VGND sg13g2_fill_1
X_5059__72 VPWR VGND net72 sg13g2_tiehi
X_4007_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\] net557 _1675_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_37_161 VPWR VGND sg13g2_decap_4
XFILLER_26_846 VPWR VGND sg13g2_decap_8
XFILLER_38_1007 VPWR VGND sg13g2_decap_8
XFILLER_25_378 VPWR VGND sg13g2_fill_1
X_4909_ net32 VGND VPWR _0337_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\]
+ net635 sg13g2_dfrbpq_1
XFILLER_5_739 VPWR VGND sg13g2_decap_8
XFILLER_1_956 VPWR VGND sg13g2_decap_8
XFILLER_49_938 VPWR VGND sg13g2_decap_8
Xhold30 serialize.n417\[6\] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold41 serialize.n410 VPWR VGND net446 sg13g2_dlygate4sd3_1
XFILLER_45_73 VPWR VGND sg13g2_fill_2
XFILLER_43_120 VPWR VGND sg13g2_fill_2
XFILLER_16_389 VPWR VGND sg13g2_fill_1
XFILLER_31_337 VPWR VGND sg13g2_fill_1
XFILLER_4_761 VPWR VGND sg13g2_decap_8
XFILLER_4_794 VPWR VGND sg13g2_decap_8
X_3240_ _0943_ _0949_ _0950_ _0321_ VPWR VGND sg13g2_nor3_1
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_3171_ _0900_ _0895_ _0897_ _0892_ _0884_ VPWR VGND sg13g2_a22oi_1
XFILLER_19_183 VPWR VGND sg13g2_fill_2
X_5027__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_35_610 VPWR VGND sg13g2_fill_2
XFILLER_35_621 VPWR VGND sg13g2_fill_1
XFILLER_22_315 VPWR VGND sg13g2_fill_2
XFILLER_23_827 VPWR VGND sg13g2_decap_8
X_2955_ _0719_ _0737_ _0792_ VPWR VGND sg13g2_nor2_2
X_2886_ _0775_ _0711_ _0771_ VPWR VGND sg13g2_nand2_2
X_4625_ net663 net713 _0055_ VPWR VGND sg13g2_nor2_1
X_4556_ VPWR _2185_ _2184_ VGND sg13g2_inv_1
X_3507_ VGND VPWR _1172_ _1174_ _1176_ _1175_ sg13g2_a21oi_1
X_4487_ _2120_ _0654_ _2119_ VPWR VGND sg13g2_xnor2_1
X_3438_ _1103_ _1101_ _1105_ _1107_ VPWR VGND sg13g2_a21o_1
X_3369_ _1047_ videogen.fancy_shader.video_y\[6\] _1046_ VPWR VGND sg13g2_xnor2_1
X_5108_ net256 VGND VPWR _0532_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\]
+ _0180_ sg13g2_dfrbpq_1
XFILLER_45_407 VPWR VGND sg13g2_fill_1
X_5039_ net166 VGND VPWR _0467_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\]
+ _0124_ sg13g2_dfrbpq_1
XFILLER_26_610 VPWR VGND sg13g2_decap_8
XFILLER_41_624 VPWR VGND sg13g2_decap_4
XFILLER_25_164 VPWR VGND sg13g2_decap_8
XFILLER_40_156 VPWR VGND sg13g2_fill_2
XFILLER_40_145 VPWR VGND sg13g2_decap_8
Xclkbuf_3_5__f_clk_regs clknet_0_clk_regs clknet_3_5__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_5191__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_21_392 VPWR VGND sg13g2_fill_2
XFILLER_31_31 VPWR VGND sg13g2_decap_8
Xoutput7 net7 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_731 VPWR VGND sg13g2_decap_8
XFILLER_1_753 VPWR VGND sg13g2_decap_8
XFILLER_49_713 VPWR VGND sg13g2_fill_1
X_5163__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_45_963 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_fill_2
XFILLER_32_646 VPWR VGND sg13g2_decap_8
XFILLER_31_145 VPWR VGND sg13g2_decap_8
XFILLER_31_167 VPWR VGND sg13g2_fill_1
X_2740_ VGND VPWR _0737_ _0710_ net585 sg13g2_or2_1
XFILLER_12_381 VPWR VGND sg13g2_fill_1
XFILLER_9_875 VPWR VGND sg13g2_decap_8
X_2671_ _0716_ _0685_ _0715_ VPWR VGND sg13g2_nand2_2
X_4410_ _0906_ VPWR _2054_ VGND _2047_ _2053_ sg13g2_o21ai_1
X_4341_ net606 VPWR _1992_ VGND tmds_green.n126 _0860_ sg13g2_o21ai_1
XFILLER_28_1006 VPWR VGND sg13g2_decap_8
X_4272_ _1899_ _1912_ _1873_ _1934_ VPWR VGND _1913_ sg13g2_nand4_1
X_3223_ VGND VPWR _0675_ _0937_ _0317_ net745 sg13g2_a21oi_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_3154_ _0882_ net547 _0883_ VPWR VGND sg13g2_xor2_1
X_3085_ net443 blue_tmds_par\[2\] net700 serialize.n429\[4\] VPWR VGND sg13g2_mux2_1
X_4890__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_35_462 VPWR VGND sg13g2_decap_4
XFILLER_35_473 VPWR VGND sg13g2_decap_8
X_3987_ net617 _1649_ _1654_ _1655_ VPWR VGND sg13g2_nor3_1
X_5198__82 VPWR VGND net82 sg13g2_tiehi
X_2938_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\] _0786_ _0400_
+ VPWR VGND sg13g2_mux2_1
X_2869_ VGND VPWR _0633_ _0768_ _0452_ _0769_ sg13g2_a21oi_1
X_4608_ net655 net707 _0038_ VPWR VGND sg13g2_nor2_1
X_4539_ VPWR _2168_ _2167_ VGND sg13g2_inv_1
XFILLER_27_963 VPWR VGND sg13g2_decap_8
XFILLER_26_473 VPWR VGND sg13g2_decap_4
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_26_495 VPWR VGND sg13g2_fill_2
XFILLER_9_105 VPWR VGND sg13g2_decap_4
XFILLER_6_834 VPWR VGND sg13g2_fill_1
XFILLER_5_344 VPWR VGND sg13g2_decap_8
XFILLER_5_399 VPWR VGND sg13g2_decap_8
XFILLER_1_550 VPWR VGND sg13g2_decap_8
XFILLER_49_576 VPWR VGND sg13g2_decap_8
XFILLER_36_226 VPWR VGND sg13g2_fill_1
XFILLER_17_440 VPWR VGND sg13g2_decap_8
XFILLER_17_451 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_fill_1
XFILLER_18_996 VPWR VGND sg13g2_decap_8
XFILLER_44_270 VPWR VGND sg13g2_decap_4
X_4890_ net70 VGND VPWR _0318_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\]
+ net631 sg13g2_dfrbpq_1
X_3910_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\] net558 _1579_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_410 VPWR VGND sg13g2_fill_1
X_3841_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\] net554 _1510_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_605 VPWR VGND sg13g2_decap_4
XFILLER_33_966 VPWR VGND sg13g2_decap_8
XFILLER_20_627 VPWR VGND sg13g2_decap_8
X_3772_ _1441_ net593 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
X_2723_ net546 _0718_ _0732_ VPWR VGND sg13g2_and2_1
X_2654_ _0705_ _0706_ net619 _0707_ VPWR VGND sg13g2_nand3_1
X_2585_ VPWR _0641_ videogen.fancy_shader.n646\[9\] VGND sg13g2_inv_1
X_4324_ _1981_ tmds_red.n102 _0914_ VPWR VGND sg13g2_xnor2_1
X_4255_ _1894_ VPWR _1917_ VGND _1877_ _1898_ sg13g2_o21ai_1
XFILLER_41_1014 VPWR VGND sg13g2_decap_8
X_3206_ _0927_ net797 _0926_ VPWR VGND sg13g2_nand2_1
X_4186_ _1836_ _1837_ _1848_ VPWR VGND _1827_ sg13g2_nand3b_1
X_3137_ tmds_red.dc_balancing_reg\[1\] tmds_red.dc_balancing_reg\[0\] tmds_red.dc_balancing_reg\[3\]
+ tmds_red.dc_balancing_reg\[2\] _0866_ VPWR VGND sg13g2_nor4_1
XFILLER_27_259 VPWR VGND sg13g2_fill_1
XFILLER_43_719 VPWR VGND sg13g2_fill_2
X_3068_ _0836_ _0849_ net7 VPWR VGND sg13g2_nor2_1
XFILLER_42_229 VPWR VGND sg13g2_fill_1
XFILLER_36_793 VPWR VGND sg13g2_decap_8
XFILLER_24_955 VPWR VGND sg13g2_decap_8
XFILLER_23_454 VPWR VGND sg13g2_decap_8
XFILLER_23_476 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_4
XFILLER_10_148 VPWR VGND sg13g2_fill_2
XFILLER_10_159 VPWR VGND sg13g2_fill_1
XFILLER_3_815 VPWR VGND sg13g2_decap_8
XFILLER_2_336 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_fill_1
Xfanout651 net654 net651 VPWR VGND sg13g2_buf_2
Xfanout640 net648 net640 VPWR VGND sg13g2_buf_8
Xfanout684 net685 net684 VPWR VGND sg13g2_buf_8
Xfanout673 net674 net673 VPWR VGND sg13g2_buf_8
Xfanout662 net672 net662 VPWR VGND sg13g2_buf_8
Xfanout695 net700 net695 VPWR VGND sg13g2_buf_8
XFILLER_42_730 VPWR VGND sg13g2_decap_8
XFILLER_15_933 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_fill_2
XFILLER_41_295 VPWR VGND sg13g2_decap_8
X_5177__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_6_642 VPWR VGND sg13g2_fill_2
XFILLER_6_697 VPWR VGND sg13g2_decap_4
XFILLER_5_141 VPWR VGND sg13g2_fill_1
X_4040_ VPWR _1705_ _1704_ VGND sg13g2_inv_1
XFILLER_37_513 VPWR VGND sg13g2_fill_1
X_4942_ net342 VGND VPWR _0370_ hsync net639 sg13g2_dfrbpq_2
XFILLER_24_229 VPWR VGND sg13g2_decap_8
XFILLER_17_292 VPWR VGND sg13g2_fill_2
XFILLER_32_240 VPWR VGND sg13g2_decap_8
X_4873_ net95 VGND VPWR _0301_ videogen.fancy_shader.video_x\[2\] net647 sg13g2_dfrbpq_2
XFILLER_20_424 VPWR VGND sg13g2_fill_1
XFILLER_21_936 VPWR VGND sg13g2_decap_8
XFILLER_32_251 VPWR VGND sg13g2_fill_1
XFILLER_20_435 VPWR VGND sg13g2_decap_4
X_3824_ _1492_ VPWR _1493_ VGND _1458_ _1468_ sg13g2_o21ai_1
X_3755_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\] net584 _1424_ VPWR
+ VGND sg13g2_nor2_1
X_2706_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\] net792 _0727_ _0582_
+ VPWR VGND sg13g2_mux2_1
X_3686_ net597 VPWR _1355_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\]
+ net580 sg13g2_o21ai_1
XFILLER_9_491 VPWR VGND sg13g2_decap_4
X_2637_ _0690_ net615 _0688_ VPWR VGND sg13g2_xnor2_1
X_4307_ _1953_ _1948_ _1950_ _1969_ VPWR VGND sg13g2_mux2_1
X_4238_ _1900_ _1877_ _1898_ VPWR VGND sg13g2_xnor2_1
X_4169_ _1820_ _1821_ _1826_ _1831_ VPWR VGND sg13g2_nor3_1
XFILLER_24_730 VPWR VGND sg13g2_decap_8
XFILLER_12_947 VPWR VGND sg13g2_decap_8
XFILLER_23_273 VPWR VGND sg13g2_fill_2
XFILLER_11_435 VPWR VGND sg13g2_decap_8
X_4920__382 VPWR VGND net382 sg13g2_tiehi
XFILLER_23_284 VPWR VGND sg13g2_fill_1
XFILLER_7_439 VPWR VGND sg13g2_decap_4
X_5090__353 VPWR VGND net353 sg13g2_tiehi
XFILLER_47_833 VPWR VGND sg13g2_fill_1
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_19_524 VPWR VGND sg13g2_fill_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_34_527 VPWR VGND sg13g2_decap_8
XFILLER_15_752 VPWR VGND sg13g2_fill_2
XFILLER_9_45 VPWR VGND sg13g2_fill_2
XFILLER_15_785 VPWR VGND sg13g2_decap_4
XFILLER_30_755 VPWR VGND sg13g2_fill_1
XFILLER_7_962 VPWR VGND sg13g2_decap_8
XFILLER_11_980 VPWR VGND sg13g2_decap_8
X_3540_ VPWR VGND _1206_ _1189_ _1201_ _1193_ _1209_ _1194_ sg13g2_a221oi_1
X_5210_ net802 VGND VPWR serialize.n428\[2\] serialize.n414\[0\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3471_ _1120_ VPWR _1140_ VGND _1116_ _1117_ sg13g2_o21ai_1
X_5141_ net69 VGND VPWR _0565_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\]
+ _0213_ sg13g2_dfrbpq_1
XFILLER_36_2 VPWR VGND sg13g2_fill_1
X_5072_ net35 VGND VPWR _0496_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\]
+ _0153_ sg13g2_dfrbpq_1
X_4023_ _1690_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1691_ VPWR VGND
+ sg13g2_nor2b_1
XFILLER_49_192 VPWR VGND sg13g2_decap_8
XFILLER_38_855 VPWR VGND sg13g2_fill_1
XFILLER_38_888 VPWR VGND sg13g2_fill_2
XFILLER_25_516 VPWR VGND sg13g2_fill_1
XFILLER_37_398 VPWR VGND sg13g2_fill_1
XFILLER_25_527 VPWR VGND sg13g2_decap_8
X_4925_ net372 VGND VPWR _0353_ videogen.fancy_shader.n646\[7\] net634 sg13g2_dfrbpq_2
XFILLER_33_571 VPWR VGND sg13g2_fill_2
X_4856_ net127 VGND VPWR _0284_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\]
+ _0015_ sg13g2_dfrbpq_1
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_21_744 VPWR VGND sg13g2_decap_4
X_3807_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\] net556 _1476_ VPWR
+ VGND sg13g2_nor2_1
X_5037__170 VPWR VGND net170 sg13g2_tiehi
X_4787_ net657 net709 _0217_ VPWR VGND sg13g2_nor2_1
X_3738_ _1407_ net594 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_4_409 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_25 VPWR VGND uio_oe[6] sg13g2_tielo
X_3669_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\] net561 _1338_ VPWR
+ VGND sg13g2_nor2_1
X_4903__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_0_648 VPWR VGND sg13g2_decap_8
XFILLER_29_844 VPWR VGND sg13g2_decap_8
XFILLER_16_516 VPWR VGND sg13g2_fill_2
XFILLER_28_354 VPWR VGND sg13g2_fill_1
XFILLER_44_858 VPWR VGND sg13g2_decap_4
XFILLER_43_335 VPWR VGND sg13g2_decap_8
XFILLER_43_324 VPWR VGND sg13g2_decap_4
XFILLER_43_313 VPWR VGND sg13g2_decap_4
X_5194__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_34_53 VPWR VGND sg13g2_decap_4
XFILLER_12_755 VPWR VGND sg13g2_decap_8
XFILLER_34_86 VPWR VGND sg13g2_fill_1
XFILLER_34_97 VPWR VGND sg13g2_decap_8
XFILLER_11_243 VPWR VGND sg13g2_decap_4
XFILLER_7_247 VPWR VGND sg13g2_decap_8
XFILLER_4_932 VPWR VGND sg13g2_decap_8
XFILLER_3_475 VPWR VGND sg13g2_decap_8
XFILLER_22_8 VPWR VGND sg13g2_decap_4
X_5068__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_34_324 VPWR VGND sg13g2_decap_8
XFILLER_22_519 VPWR VGND sg13g2_decap_4
X_2971_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\] _0795_ _0312_
+ VPWR VGND sg13g2_mux2_1
X_4710_ net679 net731 _0140_ VPWR VGND sg13g2_nor2_1
X_4641_ net664 net716 _0071_ VPWR VGND sg13g2_nor2_1
X_4572_ VGND VPWR _2198_ _2199_ _2200_ _2057_ sg13g2_a21oi_1
XFILLER_7_770 VPWR VGND sg13g2_fill_1
XFILLER_7_781 VPWR VGND sg13g2_fill_1
X_3523_ _1192_ _1190_ _1191_ VPWR VGND sg13g2_xnor2_1
X_3454_ VGND VPWR _0642_ _0651_ _1123_ _1119_ sg13g2_a21oi_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_3385_ net795 VPWR _1056_ VGND videogen.test_lut_thingy.gol_counter_reg\[3\] _1055_
+ sg13g2_o21ai_1
X_5124_ net193 VGND VPWR _0548_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\]
+ _0196_ sg13g2_dfrbpq_1
X_5055_ net98 VGND VPWR _0483_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\]
+ _0140_ sg13g2_dfrbpq_1
X_4006_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\] net588 _1674_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_26_825 VPWR VGND sg13g2_decap_8
XFILLER_25_335 VPWR VGND sg13g2_decap_8
XFILLER_25_346 VPWR VGND sg13g2_fill_1
XFILLER_13_519 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk_regs clknet_0_clk_regs clknet_3_4__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_4908_ net34 VGND VPWR _0336_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\]
+ net635 sg13g2_dfrbpq_2
XFILLER_21_563 VPWR VGND sg13g2_decap_4
X_4839_ net153 VGND VPWR _0267_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\]
+ _0006_ sg13g2_dfrbpq_1
XFILLER_21_585 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_935 VPWR VGND sg13g2_decap_8
XFILLER_49_917 VPWR VGND sg13g2_decap_8
Xhold20 serialize.n417\[7\] VPWR VGND net425 sg13g2_dlygate4sd3_1
XFILLER_48_416 VPWR VGND sg13g2_fill_2
Xhold31 serialize.n414\[2\] VPWR VGND net436 sg13g2_dlygate4sd3_1
XFILLER_0_467 VPWR VGND sg13g2_decap_8
XFILLER_17_836 VPWR VGND sg13g2_decap_4
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_16_368 VPWR VGND sg13g2_fill_1
XFILLER_40_894 VPWR VGND sg13g2_decap_8
XFILLER_40_883 VPWR VGND sg13g2_decap_4
XFILLER_8_534 VPWR VGND sg13g2_decap_8
XFILLER_12_596 VPWR VGND sg13g2_fill_2
XFILLER_6_24 VPWR VGND sg13g2_decap_8
XFILLER_6_13 VPWR VGND sg13g2_fill_2
X_3170_ _0899_ _0898_ _0888_ VPWR VGND sg13g2_nand2b_1
XFILLER_13_4 VPWR VGND sg13g2_decap_4
XFILLER_23_806 VPWR VGND sg13g2_fill_2
X_2954_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\] _0791_ _0389_
+ VPWR VGND sg13g2_mux2_1
X_2885_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\] net784 _0774_ _0441_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_371 VPWR VGND sg13g2_decap_8
XFILLER_30_382 VPWR VGND sg13g2_fill_1
X_5151__320 VPWR VGND net320 sg13g2_tiehi
X_4624_ net663 net715 _0054_ VPWR VGND sg13g2_nor2_1
X_4555_ _2148_ _2181_ _2184_ VPWR VGND sg13g2_nor2_1
X_3506_ _1149_ _1168_ _1175_ VPWR VGND sg13g2_and2_1
X_4486_ VGND VPWR tmds_green.dc_balancing_reg\[3\] _2086_ _2119_ _2084_ sg13g2_a21oi_1
X_3437_ VGND VPWR _1101_ _1103_ _1106_ _1105_ sg13g2_a21oi_1
X_4885__79 VPWR VGND net79 sg13g2_tiehi
X_3368_ net745 _1045_ _1046_ _0361_ VPWR VGND sg13g2_nor3_1
X_5107_ net260 VGND VPWR _0531_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\]
+ _0179_ sg13g2_dfrbpq_1
XFILLER_46_909 VPWR VGND sg13g2_decap_8
X_3299_ _0985_ VPWR _0991_ VGND _0986_ _0988_ sg13g2_o21ai_1
XFILLER_39_983 VPWR VGND sg13g2_decap_8
X_5038_ net168 VGND VPWR _0466_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\]
+ _0123_ sg13g2_dfrbpq_1
XFILLER_5_504 VPWR VGND sg13g2_fill_2
Xoutput8 net8 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_0_220 VPWR VGND sg13g2_decap_8
XFILLER_0_253 VPWR VGND sg13g2_decap_8
XFILLER_48_202 VPWR VGND sg13g2_decap_8
XFILLER_36_408 VPWR VGND sg13g2_decap_4
XFILLER_36_419 VPWR VGND sg13g2_fill_1
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_16_132 VPWR VGND sg13g2_decap_8
XFILLER_17_633 VPWR VGND sg13g2_fill_2
XFILLER_44_474 VPWR VGND sg13g2_fill_1
XFILLER_16_187 VPWR VGND sg13g2_decap_4
XFILLER_31_124 VPWR VGND sg13g2_decap_8
XFILLER_32_625 VPWR VGND sg13g2_fill_2
XFILLER_9_832 VPWR VGND sg13g2_decap_8
XFILLER_13_883 VPWR VGND sg13g2_fill_2
XFILLER_8_364 VPWR VGND sg13g2_fill_1
XFILLER_8_342 VPWR VGND sg13g2_decap_8
X_2670_ _0715_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] _0688_ VPWR VGND
+ sg13g2_nand2_1
X_4340_ VGND VPWR _0654_ net606 _0505_ net748 sg13g2_a21oi_1
X_4271_ _1932_ VPWR _1933_ VGND _1903_ _1910_ sg13g2_o21ai_1
X_3222_ _0935_ _0936_ _0937_ VPWR VGND sg13g2_nor2_1
X_3153_ _0882_ tmds_red.n100 tmds_red.n102 VPWR VGND sg13g2_xnor2_1
X_3084_ net433 blue_tmds_par\[3\] net700 serialize.n429\[3\] VPWR VGND sg13g2_mux2_1
XFILLER_36_920 VPWR VGND sg13g2_decap_4
XFILLER_47_290 VPWR VGND sg13g2_fill_1
XFILLER_35_430 VPWR VGND sg13g2_decap_8
XFILLER_36_997 VPWR VGND sg13g2_decap_8
XFILLER_23_647 VPWR VGND sg13g2_decap_8
X_3986_ net625 _1650_ _1651_ _1653_ _1654_ VPWR VGND sg13g2_nor4_1
XFILLER_23_658 VPWR VGND sg13g2_decap_8
X_2937_ _0786_ _0781_ VPWR VGND _0726_ sg13g2_nand2b_2
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
X_2868_ net757 _0768_ _0769_ VPWR VGND sg13g2_nor2_1
X_4607_ net683 net719 _0037_ VPWR VGND sg13g2_nor2_1
X_2799_ _0700_ _0728_ _0752_ VPWR VGND sg13g2_nor2_2
X_4538_ _2167_ _2141_ _2166_ VPWR VGND sg13g2_nand2_1
Xfanout800 net801 net800 VPWR VGND sg13g2_buf_2
X_4469_ _2085_ net600 _2089_ _2103_ VPWR VGND sg13g2_a21o_1
XFILLER_46_706 VPWR VGND sg13g2_fill_1
XFILLER_19_909 VPWR VGND sg13g2_decap_8
XFILLER_27_942 VPWR VGND sg13g2_decap_8
XFILLER_26_43 VPWR VGND sg13g2_fill_1
XFILLER_26_65 VPWR VGND sg13g2_decap_8
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_5_334 VPWR VGND sg13g2_decap_4
X_4930__362 VPWR VGND net362 sg13g2_tiehi
XFILLER_3_58 VPWR VGND sg13g2_decap_8
XFILLER_49_555 VPWR VGND sg13g2_decap_8
XFILLER_37_706 VPWR VGND sg13g2_fill_1
XFILLER_18_975 VPWR VGND sg13g2_decap_8
XFILLER_33_945 VPWR VGND sg13g2_decap_8
X_3840_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\] net576 _1509_ VPWR
+ VGND sg13g2_nor2_1
X_3771_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\] net563 _1440_ VPWR
+ VGND sg13g2_nor2_1
X_2722_ net792 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\] _0731_ _0570_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_651 VPWR VGND sg13g2_fill_2
XFILLER_8_150 VPWR VGND sg13g2_fill_1
XFILLER_9_684 VPWR VGND sg13g2_fill_1
XFILLER_8_194 VPWR VGND sg13g2_decap_8
X_2653_ _0647_ net595 _0684_ _0706_ VPWR VGND sg13g2_nor3_1
X_2584_ VPWR _0640_ videogen.fancy_shader.video_y\[2\] VGND sg13g2_inv_1
X_4323_ _1980_ VPWR _0383_ VGND net748 _1976_ sg13g2_o21ai_1
X_4254_ _1916_ _1913_ _1915_ VPWR VGND sg13g2_nand2_1
X_3205_ _0926_ _0813_ videogen.fancy_shader.video_x\[4\] VPWR VGND sg13g2_nand2b_1
X_4185_ VPWR _1847_ _1846_ VGND sg13g2_inv_1
X_3136_ VGND VPWR _0861_ _0864_ _0273_ _0865_ sg13g2_a21oi_1
X_3067_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\] _0846_ _0849_
+ _0848_ sg13g2_a21oi_1
XFILLER_24_934 VPWR VGND sg13g2_decap_8
XFILLER_35_293 VPWR VGND sg13g2_fill_1
XFILLER_12_12 VPWR VGND sg13g2_decap_8
X_3969_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\] net575 _1637_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_2_359 VPWR VGND sg13g2_decap_8
Xfanout630 net631 net630 VPWR VGND sg13g2_buf_8
Xfanout641 net643 net641 VPWR VGND sg13g2_buf_8
Xfanout663 net666 net663 VPWR VGND sg13g2_buf_8
Xfanout685 net687 net685 VPWR VGND sg13g2_buf_8
Xfanout674 net682 net674 VPWR VGND sg13g2_buf_8
Xfanout652 net653 net652 VPWR VGND sg13g2_buf_8
Xfanout696 net699 net696 VPWR VGND sg13g2_buf_8
XFILLER_37_20 VPWR VGND sg13g2_fill_1
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
XFILLER_15_912 VPWR VGND sg13g2_decap_8
XFILLER_33_208 VPWR VGND sg13g2_fill_2
XFILLER_15_989 VPWR VGND sg13g2_decap_8
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_fill_2
XFILLER_1_370 VPWR VGND sg13g2_fill_1
XFILLER_49_330 VPWR VGND sg13g2_decap_4
XFILLER_49_352 VPWR VGND sg13g2_decap_4
X_4941_ net343 VGND VPWR _0369_ videogen.test_lut_thingy.gol_counter_reg\[3\] net639
+ sg13g2_dfrbpq_1
X_4872_ net96 VGND VPWR _0300_ videogen.fancy_shader.video_x\[1\] net647 sg13g2_dfrbpq_2
XFILLER_21_915 VPWR VGND sg13g2_decap_8
X_3823_ _1491_ net610 _1492_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_263 VPWR VGND sg13g2_fill_2
XFILLER_32_274 VPWR VGND sg13g2_decap_8
XFILLER_20_458 VPWR VGND sg13g2_decap_8
X_3754_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\] net561 _1423_ VPWR
+ VGND sg13g2_nor2_1
X_2705_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\] net782 _0727_ _0583_
+ VPWR VGND sg13g2_mux2_1
X_3685_ _1350_ _1351_ _1352_ _1353_ _1354_ VPWR VGND sg13g2_nor4_1
X_2636_ net614 net620 net585 _0689_ VPWR VGND sg13g2_nor3_1
X_4306_ _1968_ _1949_ _1955_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_90 VPWR VGND sg13g2_fill_2
X_4237_ _1898_ _1877_ _1899_ VPWR VGND sg13g2_xor2_1
XFILLER_28_503 VPWR VGND sg13g2_decap_8
X_4168_ _1829_ _1828_ _1830_ VPWR VGND sg13g2_xor2_1
X_3119_ tmds_green.dc_balancing_reg\[0\] _0852_ _0263_ VPWR VGND sg13g2_and2_1
X_4099_ VGND VPWR _1747_ _1752_ _1764_ _1750_ sg13g2_a21oi_1
XFILLER_12_926 VPWR VGND sg13g2_decap_8
XFILLER_8_919 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_2_134 VPWR VGND sg13g2_decap_4
XFILLER_2_156 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_48_96 VPWR VGND sg13g2_fill_2
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_46_366 VPWR VGND sg13g2_fill_2
XFILLER_46_355 VPWR VGND sg13g2_fill_1
XFILLER_0_48 VPWR VGND sg13g2_fill_2
XFILLER_19_569 VPWR VGND sg13g2_fill_2
XFILLER_46_377 VPWR VGND sg13g2_fill_2
XFILLER_15_797 VPWR VGND sg13g2_decap_8
XFILLER_30_723 VPWR VGND sg13g2_decap_4
XFILLER_7_941 VPWR VGND sg13g2_decap_8
X_3470_ _1134_ _1136_ _1139_ VPWR VGND sg13g2_nor2_2
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_5140_ net78 VGND VPWR _0564_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\]
+ _0212_ sg13g2_dfrbpq_1
X_5071_ net39 VGND VPWR _0495_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\]
+ _0152_ sg13g2_dfrbpq_1
X_4022_ net611 _1678_ _1689_ _1690_ VPWR VGND sg13g2_nor3_1
XFILLER_49_171 VPWR VGND sg13g2_decap_8
XFILLER_37_333 VPWR VGND sg13g2_fill_2
X_5182__293 VPWR VGND net293 sg13g2_tiehi
XFILLER_38_867 VPWR VGND sg13g2_decap_8
XFILLER_37_355 VPWR VGND sg13g2_decap_4
Xclkbuf_3_3__f_clk_regs clknet_0_clk_regs clknet_3_3__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_4924_ net374 VGND VPWR _0352_ videogen.fancy_shader.n646\[6\] net634 sg13g2_dfrbpq_2
XFILLER_21_701 VPWR VGND sg13g2_decap_8
X_4855_ net129 VGND VPWR _0283_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\]
+ _0014_ sg13g2_dfrbpq_1
X_4786_ net658 net710 _0216_ VPWR VGND sg13g2_nor2_1
X_3806_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\] net588 _1475_ VPWR
+ VGND sg13g2_nor2_1
X_3737_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\] net569 _1406_ VPWR
+ VGND sg13g2_nor2_1
X_3668_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\] net551 _1337_ VPWR
+ VGND sg13g2_nor2_1
Xheichips25_bagel_26 VPWR VGND uio_oe[7] sg13g2_tielo
X_2619_ _0672_ VPWR _0262_ VGND net415 serialize.n433\[1\] sg13g2_o21ai_1
X_3599_ VPWR _1268_ _1267_ VGND sg13g2_inv_1
XFILLER_0_616 VPWR VGND sg13g2_decap_4
XFILLER_18_44 VPWR VGND sg13g2_fill_2
XFILLER_12_712 VPWR VGND sg13g2_fill_1
XFILLER_34_32 VPWR VGND sg13g2_fill_1
XFILLER_11_288 VPWR VGND sg13g2_fill_1
XFILLER_11_299 VPWR VGND sg13g2_decap_8
XFILLER_4_911 VPWR VGND sg13g2_decap_8
XFILLER_4_988 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_38_108 VPWR VGND sg13g2_decap_8
XFILLER_47_620 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_decap_8
XFILLER_46_185 VPWR VGND sg13g2_decap_4
XFILLER_46_174 VPWR VGND sg13g2_fill_1
XFILLER_15_550 VPWR VGND sg13g2_decap_4
X_2970_ _0795_ _0720_ VPWR VGND _0714_ sg13g2_nand2b_2
X_4640_ net664 net715 _0070_ VPWR VGND sg13g2_nor2_1
X_4571_ _2189_ _2061_ _2199_ VPWR VGND _2175_ sg13g2_nand3b_1
X_3522_ VGND VPWR _0991_ _0993_ _1191_ _0992_ sg13g2_a21oi_1
X_3453_ _1121_ VPWR _1122_ VGND _1116_ _1117_ sg13g2_o21ai_1
X_3384_ net751 _1054_ _1055_ _0368_ VPWR VGND sg13g2_nor3_1
X_5123_ net197 VGND VPWR _0547_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\]
+ _0195_ sg13g2_dfrbpq_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_29_108 VPWR VGND sg13g2_decap_8
X_5054_ net102 VGND VPWR _0482_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\]
+ _0139_ sg13g2_dfrbpq_1
X_4005_ net624 VPWR _1673_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\]
+ net570 sg13g2_o21ai_1
XFILLER_26_804 VPWR VGND sg13g2_decap_8
X_5080__375 VPWR VGND net375 sg13g2_tiehi
XFILLER_25_358 VPWR VGND sg13g2_fill_1
XFILLER_25_369 VPWR VGND sg13g2_decap_8
X_4907_ net36 VGND VPWR _0335_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ net635 sg13g2_dfrbpq_1
X_4838_ net154 VGND VPWR net743 clockdiv.q2temp net405 sg13g2_dfrbpq_1
X_4769_ net683 net734 _0199_ VPWR VGND sg13g2_nor2_1
XFILLER_1_914 VPWR VGND sg13g2_decap_8
XFILLER_0_446 VPWR VGND sg13g2_decap_8
Xhold32 serialize.n417\[2\] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xhold10 _0004_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold21 serialize.n411\[5\] VPWR VGND net426 sg13g2_dlygate4sd3_1
XFILLER_29_76 VPWR VGND sg13g2_decap_8
XFILLER_21_1013 VPWR VGND sg13g2_decap_8
XFILLER_29_664 VPWR VGND sg13g2_fill_2
XFILLER_44_623 VPWR VGND sg13g2_fill_1
XFILLER_16_314 VPWR VGND sg13g2_fill_2
XFILLER_43_122 VPWR VGND sg13g2_fill_1
XFILLER_28_185 VPWR VGND sg13g2_fill_2
XFILLER_45_86 VPWR VGND sg13g2_fill_2
XFILLER_45_75 VPWR VGND sg13g2_fill_1
X_4957__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_8_579 VPWR VGND sg13g2_fill_1
XFILLER_4_730 VPWR VGND sg13g2_decap_8
XFILLER_3_273 VPWR VGND sg13g2_decap_8
XFILLER_48_984 VPWR VGND sg13g2_decap_8
XFILLER_16_870 VPWR VGND sg13g2_fill_1
XFILLER_22_339 VPWR VGND sg13g2_decap_4
XFILLER_34_177 VPWR VGND sg13g2_decap_4
X_2953_ net776 videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\] _0791_ _0390_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_851 VPWR VGND sg13g2_fill_2
X_2884_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\] net773 _0774_ _0442_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_350 VPWR VGND sg13g2_fill_2
X_4623_ net661 net713 _0053_ VPWR VGND sg13g2_nor2_1
X_4554_ VGND VPWR net602 _2175_ _2183_ _2182_ sg13g2_a21oi_1
XFILLER_7_590 VPWR VGND sg13g2_fill_1
X_3505_ VGND VPWR _1149_ _1158_ _1174_ _1167_ sg13g2_a21oi_1
X_4485_ _2106_ VPWR _2118_ VGND _2101_ _2103_ sg13g2_o21ai_1
XFILLER_44_1013 VPWR VGND sg13g2_decap_8
X_3436_ _1105_ videogen.fancy_shader.video_y\[8\] net609 VPWR VGND sg13g2_xnor2_1
X_3367_ videogen.fancy_shader.video_y\[5\] _1044_ _1046_ VPWR VGND sg13g2_and2_1
X_5106_ net268 VGND VPWR _0530_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\]
+ _0178_ sg13g2_dfrbpq_1
X_5037_ net170 VGND VPWR _0465_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\]
+ _0122_ sg13g2_dfrbpq_1
X_3298_ _0990_ _0987_ _0989_ VPWR VGND sg13g2_nand2_2
X_5006__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_38_461 VPWR VGND sg13g2_fill_1
XFILLER_38_450 VPWR VGND sg13g2_decap_4
XFILLER_13_317 VPWR VGND sg13g2_fill_1
XFILLER_13_328 VPWR VGND sg13g2_decap_4
XFILLER_15_45 VPWR VGND sg13g2_decap_4
XFILLER_22_862 VPWR VGND sg13g2_decap_8
XFILLER_31_11 VPWR VGND sg13g2_fill_2
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_5_549 VPWR VGND sg13g2_fill_2
X_4917__388 VPWR VGND net388 sg13g2_tiehi
XFILLER_1_700 VPWR VGND sg13g2_decap_8
Xoutput11 net11 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_out[3] VPWR VGND sg13g2_buf_1
X_5087__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_1_788 VPWR VGND sg13g2_decap_8
XFILLER_45_921 VPWR VGND sg13g2_decap_8
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_16_155 VPWR VGND sg13g2_decap_8
XFILLER_16_177 VPWR VGND sg13g2_fill_1
XFILLER_31_103 VPWR VGND sg13g2_decap_4
XFILLER_31_114 VPWR VGND sg13g2_fill_1
XFILLER_13_862 VPWR VGND sg13g2_decap_8
XFILLER_8_376 VPWR VGND sg13g2_fill_2
X_4853__133 VPWR VGND net133 sg13g2_tiehi
X_4270_ _1900_ VPWR _1932_ VGND _1902_ _1910_ sg13g2_o21ai_1
X_5146__401 VPWR VGND net401 sg13g2_tiehi
X_3221_ _0936_ videogen.fancy_shader.video_y\[1\] net608 VPWR VGND sg13g2_xnor2_1
XFILLER_39_225 VPWR VGND sg13g2_fill_2
X_3152_ VGND VPWR tmds_red.n100 _0880_ _0881_ _0878_ sg13g2_a21oi_1
X_3083_ net437 blue_tmds_par\[2\] net694 serialize.n429\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_36_976 VPWR VGND sg13g2_decap_8
X_3985_ _1652_ VPWR _1653_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\]
+ net558 sg13g2_o21ai_1
XFILLER_22_147 VPWR VGND sg13g2_decap_8
XFILLER_22_158 VPWR VGND sg13g2_decap_8
X_2936_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\] net784 _0785_ _0401_
+ VPWR VGND sg13g2_mux2_1
X_2867_ _0768_ _0716_ _0757_ VPWR VGND sg13g2_nand2_2
XFILLER_30_191 VPWR VGND sg13g2_fill_2
X_5201__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_31_692 VPWR VGND sg13g2_decap_8
X_4606_ net684 net736 _0036_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
X_2798_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\] net789 _0751_ _0514_
+ VPWR VGND sg13g2_mux2_1
XFILLER_2_519 VPWR VGND sg13g2_decap_8
X_4537_ _2166_ tmds_blue.n193 _2165_ VPWR VGND sg13g2_nand2_1
X_4468_ VPWR _2102_ _2101_ VGND sg13g2_inv_1
Xfanout801 net806 net801 VPWR VGND sg13g2_buf_8
X_3419_ _1086_ _1087_ _1088_ VPWR VGND sg13g2_nor2_1
X_4399_ _0910_ _2029_ _2044_ VPWR VGND _2030_ sg13g2_nand3b_1
X_4947__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_27_921 VPWR VGND sg13g2_decap_8
XFILLER_45_228 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_fill_2
XFILLER_27_998 VPWR VGND sg13g2_decap_8
XFILLER_41_401 VPWR VGND sg13g2_decap_8
XFILLER_13_114 VPWR VGND sg13g2_fill_1
XFILLER_14_615 VPWR VGND sg13g2_decap_8
XFILLER_13_125 VPWR VGND sg13g2_decap_4
XFILLER_6_803 VPWR VGND sg13g2_fill_2
XFILLER_10_843 VPWR VGND sg13g2_fill_2
XFILLER_6_814 VPWR VGND sg13g2_fill_1
XFILLER_5_324 VPWR VGND sg13g2_fill_2
XFILLER_5_357 VPWR VGND sg13g2_decap_4
XFILLER_3_26 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_fill_1
X_5167__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_18_954 VPWR VGND sg13g2_decap_8
XFILLER_29_280 VPWR VGND sg13g2_fill_2
XFILLER_45_751 VPWR VGND sg13g2_decap_4
XFILLER_32_401 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
X_3770_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\] net575 _1439_ VPWR
+ VGND sg13g2_nor2_1
X_2721_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\] _0731_ _0571_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_630 VPWR VGND sg13g2_decap_8
XFILLER_8_173 VPWR VGND sg13g2_decap_8
X_2652_ _0705_ _0685_ _0703_ VPWR VGND sg13g2_nand2_1
X_2583_ VPWR _0639_ videogen.fancy_shader.video_y\[7\] VGND sg13g2_inv_1
X_4322_ _1799_ _1979_ _1980_ VPWR VGND sg13g2_and2_1
X_4253_ _1872_ _1900_ _1915_ VPWR VGND sg13g2_nor2_1
X_3204_ _0812_ _0925_ _0302_ VPWR VGND sg13g2_nor2_1
X_4184_ _1836_ _1837_ _1846_ VPWR VGND sg13g2_and2_1
X_3135_ _0852_ VPWR _0865_ VGND _0861_ _0864_ sg13g2_o21ai_1
XFILLER_28_729 VPWR VGND sg13g2_decap_8
X_3066_ _0835_ VPWR _0848_ VGND videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ _0846_ sg13g2_o21ai_1
XFILLER_24_913 VPWR VGND sg13g2_decap_8
XFILLER_23_401 VPWR VGND sg13g2_decap_8
XFILLER_23_467 VPWR VGND sg13g2_decap_4
X_3968_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\] net563 _1636_ VPWR
+ VGND sg13g2_nor2_1
X_2919_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\] _0782_ _0415_
+ VPWR VGND sg13g2_mux2_1
X_3899_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\] net581 _1568_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_2_316 VPWR VGND sg13g2_decap_4
Xfanout631 net648 net631 VPWR VGND sg13g2_buf_8
Xfanout620 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\] net620 VPWR VGND
+ sg13g2_buf_8
Xfanout642 net643 net642 VPWR VGND sg13g2_buf_1
Xfanout664 net666 net664 VPWR VGND sg13g2_buf_2
Xfanout653 net654 net653 VPWR VGND sg13g2_buf_8
Xfanout675 net682 net675 VPWR VGND sg13g2_buf_8
Xfanout697 net699 net697 VPWR VGND sg13g2_buf_8
Xfanout686 net687 net686 VPWR VGND sg13g2_buf_1
XFILLER_37_32 VPWR VGND sg13g2_decap_8
XFILLER_18_239 VPWR VGND sg13g2_fill_2
XFILLER_42_765 VPWR VGND sg13g2_fill_2
XFILLER_15_968 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_6_611 VPWR VGND sg13g2_decap_8
XFILLER_6_600 VPWR VGND sg13g2_decap_4
XFILLER_6_644 VPWR VGND sg13g2_fill_1
XFILLER_6_688 VPWR VGND sg13g2_fill_2
XFILLER_6_677 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_fill_2
XFILLER_2_894 VPWR VGND sg13g2_decap_8
XFILLER_49_320 VPWR VGND sg13g2_fill_2
XFILLER_37_504 VPWR VGND sg13g2_decap_4
XFILLER_49_397 VPWR VGND sg13g2_decap_8
Xclkbuf_3_2__f_clk_regs clknet_0_clk_regs clknet_3_2__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_18_784 VPWR VGND sg13g2_fill_1
X_4940_ net344 VGND VPWR _0368_ videogen.test_lut_thingy.gol_counter_reg\[2\] net639
+ sg13g2_dfrbpq_1
X_4871_ net97 VGND VPWR _0299_ videogen.fancy_shader.video_x\[0\] net647 sg13g2_dfrbpq_2
X_3822_ net611 _1479_ _1490_ _1491_ VPWR VGND sg13g2_nor3_1
XFILLER_20_404 VPWR VGND sg13g2_decap_8
XFILLER_33_776 VPWR VGND sg13g2_decap_8
X_5076__391 VPWR VGND net391 sg13g2_tiehi
X_3753_ _1422_ net613 _1421_ VPWR VGND sg13g2_nand2b_1
X_3684_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\] net553 _1353_ VPWR
+ VGND sg13g2_nor2_1
X_2704_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\] net770 _0727_ _0584_
+ VPWR VGND sg13g2_mux2_1
X_2635_ net619 net587 _0688_ VPWR VGND sg13g2_nor2_1
X_4305_ VGND VPWR _1860_ _1864_ _1967_ _1857_ sg13g2_a21oi_1
XFILLER_4_80 VPWR VGND sg13g2_fill_2
X_4236_ VGND VPWR _1897_ _1898_ _1896_ _1890_ sg13g2_a21oi_2
X_4167_ _1829_ _1073_ _1706_ VPWR VGND sg13g2_xnor2_1
X_3118_ _0853_ net607 net799 VPWR VGND sg13g2_nand2_1
X_4098_ _1761_ _1760_ _1758_ _1763_ VPWR VGND sg13g2_a21o_1
XFILLER_28_559 VPWR VGND sg13g2_decap_8
X_3049_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] VPWR _0836_ VGND _0828_
+ _0835_ sg13g2_o21ai_1
XFILLER_12_905 VPWR VGND sg13g2_decap_8
XFILLER_24_765 VPWR VGND sg13g2_decap_8
XFILLER_23_275 VPWR VGND sg13g2_fill_1
XFILLER_2_113 VPWR VGND sg13g2_decap_4
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_fill_1
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_24_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_813 VPWR VGND sg13g2_decap_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_46_312 VPWR VGND sg13g2_fill_1
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_19_559 VPWR VGND sg13g2_fill_2
X_5125__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_27_592 VPWR VGND sg13g2_fill_1
XFILLER_15_765 VPWR VGND sg13g2_decap_8
XFILLER_15_776 VPWR VGND sg13g2_fill_1
XFILLER_9_47 VPWR VGND sg13g2_fill_1
XFILLER_30_735 VPWR VGND sg13g2_decap_8
XFILLER_7_920 VPWR VGND sg13g2_decap_8
XFILLER_31_1026 VPWR VGND sg13g2_fill_2
XFILLER_6_441 VPWR VGND sg13g2_fill_2
XFILLER_6_430 VPWR VGND sg13g2_decap_8
XFILLER_7_997 VPWR VGND sg13g2_decap_8
X_5070_ net43 VGND VPWR _0494_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\]
+ _0151_ sg13g2_dfrbpq_1
XFILLER_2_691 VPWR VGND sg13g2_fill_2
XFILLER_49_150 VPWR VGND sg13g2_decap_8
X_4021_ net616 _1683_ _1688_ _1689_ VPWR VGND sg13g2_nor3_1
XFILLER_38_846 VPWR VGND sg13g2_decap_8
X_4923_ net376 VGND VPWR _0351_ videogen.fancy_shader.n646\[5\] net632 sg13g2_dfrbpq_2
XFILLER_33_540 VPWR VGND sg13g2_fill_1
X_4854_ net131 VGND VPWR _0282_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\]
+ _0013_ sg13g2_dfrbpq_1
X_3805_ net624 VPWR _1474_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\]
+ net567 sg13g2_o21ai_1
X_4785_ net667 net720 _0215_ VPWR VGND sg13g2_nor2_1
X_3736_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\] net559 _1405_ VPWR
+ VGND sg13g2_nor2_1
Xheichips25_bagel_27 VPWR VGND uio_out[1] sg13g2_tielo
X_3667_ net614 VPWR _1336_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\]
+ net584 sg13g2_o21ai_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_2618_ _0672_ net415 _0671_ VPWR VGND sg13g2_nand2_1
X_3598_ _1267_ _1076_ _1265_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_628 VPWR VGND sg13g2_fill_1
X_4219_ _1881_ _1166_ _1880_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_813 VPWR VGND sg13g2_decap_8
XFILLER_28_301 VPWR VGND sg13g2_fill_1
X_5199_ net65 VGND VPWR net407 clockdiv.q0 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_29_824 VPWR VGND sg13g2_fill_2
XFILLER_16_518 VPWR VGND sg13g2_fill_1
XFILLER_28_367 VPWR VGND sg13g2_fill_2
XFILLER_12_724 VPWR VGND sg13g2_decap_8
XFILLER_12_735 VPWR VGND sg13g2_fill_1
XFILLER_34_66 VPWR VGND sg13g2_fill_2
XFILLER_11_256 VPWR VGND sg13g2_decap_8
XFILLER_7_216 VPWR VGND sg13g2_decap_4
X_5016__212 VPWR VGND net212 sg13g2_tiehi
X_5051__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_4_967 VPWR VGND sg13g2_decap_8
XFILLER_3_444 VPWR VGND sg13g2_decap_4
XFILLER_47_654 VPWR VGND sg13g2_fill_2
XFILLER_47_643 VPWR VGND sg13g2_decap_8
X_4927__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_35_838 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_fill_1
X_4973__300 VPWR VGND net300 sg13g2_tiehi
X_4570_ _2060_ VPWR _2198_ VGND _2184_ _2197_ sg13g2_o21ai_1
XFILLER_30_587 VPWR VGND sg13g2_decap_8
XFILLER_30_598 VPWR VGND sg13g2_fill_1
X_3521_ videogen.fancy_shader.n646\[3\] videogen.fancy_shader.video_y\[3\] _1190_
+ VPWR VGND sg13g2_xor2_1
X_3452_ _1118_ _1120_ _1121_ VPWR VGND sg13g2_nor2b_1
X_4897__56 VPWR VGND net56 sg13g2_tiehi
X_3383_ _1055_ videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ videogen.test_lut_thingy.gol_counter_reg\[2\] VPWR VGND sg13g2_and3_1
X_5122_ net201 VGND VPWR _0546_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\]
+ _0194_ sg13g2_dfrbpq_1
X_5053_ net106 VGND VPWR _0481_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\]
+ _0138_ sg13g2_dfrbpq_1
XFILLER_38_654 VPWR VGND sg13g2_decap_4
X_4863__113 VPWR VGND net113 sg13g2_tiehi
X_4004_ net623 _1668_ _1669_ _1671_ _1672_ VPWR VGND sg13g2_nor4_1
X_4906_ net38 VGND VPWR _0334_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\]
+ net635 sg13g2_dfrbpq_1
X_4837_ net155 VGND VPWR _0266_ clockdiv.q2 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
X_4768_ net687 net735 _0198_ VPWR VGND sg13g2_nor2_1
X_3719_ net596 VPWR _1388_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\]
+ net556 sg13g2_o21ai_1
XFILLER_4_219 VPWR VGND sg13g2_fill_2
XFILLER_4_208 VPWR VGND sg13g2_decap_8
X_4699_ net680 net730 _0129_ VPWR VGND sg13g2_nor2_1
Xhold22 serialize.n417\[5\] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold11 _0262_ VPWR VGND net416 sg13g2_dlygate4sd3_1
Xhold33 serialize.n414\[7\] VPWR VGND net438 sg13g2_dlygate4sd3_1
XFILLER_28_120 VPWR VGND sg13g2_fill_2
XFILLER_28_175 VPWR VGND sg13g2_decap_4
XFILLER_29_698 VPWR VGND sg13g2_fill_2
XFILLER_45_32 VPWR VGND sg13g2_fill_2
XFILLER_16_337 VPWR VGND sg13g2_decap_8
XFILLER_16_359 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_fill_2
XFILLER_43_178 VPWR VGND sg13g2_decap_4
XFILLER_24_370 VPWR VGND sg13g2_decap_4
XFILLER_25_893 VPWR VGND sg13g2_decap_8
XFILLER_24_392 VPWR VGND sg13g2_fill_2
XFILLER_6_15 VPWR VGND sg13g2_fill_1
X_4879__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_6_1019 VPWR VGND sg13g2_decap_4
XFILLER_0_992 VPWR VGND sg13g2_decap_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
XFILLER_47_440 VPWR VGND sg13g2_fill_2
XFILLER_37_1021 VPWR VGND sg13g2_decap_8
X_2952_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\] _0791_ _0391_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_392 VPWR VGND sg13g2_decap_8
X_2883_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\] net763 _0774_ _0443_
+ VPWR VGND sg13g2_mux2_1
X_4622_ net667 net720 _0052_ VPWR VGND sg13g2_nor2_1
X_4553_ _2057_ VPWR _2182_ VGND net602 _2181_ sg13g2_o21ai_1
X_4484_ net571 _2117_ _0621_ VPWR VGND sg13g2_nor2_1
X_3504_ _1158_ _1167_ _1173_ VPWR VGND sg13g2_nor2_2
X_3435_ net609 videogen.fancy_shader.video_y\[8\] _1104_ VPWR VGND sg13g2_xor2_1
X_3366_ videogen.fancy_shader.video_y\[5\] _1044_ _1045_ VPWR VGND sg13g2_nor2_1
X_5105_ net271 VGND VPWR _0529_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\]
+ _0177_ sg13g2_dfrbpq_1
X_3297_ videogen.fancy_shader.n646\[0\] net608 _0989_ VPWR VGND sg13g2_xor2_1
X_5036_ net172 VGND VPWR _0464_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[3\]
+ _0121_ sg13g2_dfrbpq_1
XFILLER_38_484 VPWR VGND sg13g2_fill_2
XFILLER_25_112 VPWR VGND sg13g2_fill_1
XFILLER_26_668 VPWR VGND sg13g2_fill_1
XFILLER_26_679 VPWR VGND sg13g2_decap_8
XFILLER_25_189 VPWR VGND sg13g2_decap_4
X_5062__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_5_506 VPWR VGND sg13g2_fill_1
XFILLER_31_45 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_fill_2
Xoutput12 net12 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_745 VPWR VGND sg13g2_fill_2
XFILLER_1_767 VPWR VGND sg13g2_decap_8
X_4884__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_44_432 VPWR VGND sg13g2_fill_1
XFILLER_44_421 VPWR VGND sg13g2_decap_8
XFILLER_16_112 VPWR VGND sg13g2_decap_4
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_44_487 VPWR VGND sg13g2_decap_8
XFILLER_32_627 VPWR VGND sg13g2_fill_1
XFILLER_9_801 VPWR VGND sg13g2_fill_2
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_9_812 VPWR VGND sg13g2_decap_8
XFILLER_13_885 VPWR VGND sg13g2_fill_1
XFILLER_9_889 VPWR VGND sg13g2_decap_8
X_3220_ _0935_ videogen.fancy_shader.video_y\[3\] _0640_ VPWR VGND sg13g2_nand2_1
X_3151_ _0879_ _0873_ _0880_ VPWR VGND sg13g2_xor2_1
X_3082_ net440 blue_tmds_par\[1\] net694 serialize.n429\[1\] VPWR VGND sg13g2_mux2_1
XFILLER_35_410 VPWR VGND sg13g2_fill_2
XFILLER_23_627 VPWR VGND sg13g2_fill_2
XFILLER_35_487 VPWR VGND sg13g2_decap_8
X_3984_ VGND VPWR _1652_ net568 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\]
+ sg13g2_or2_1
X_2935_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\] net773 _0785_ _0402_
+ VPWR VGND sg13g2_mux2_1
X_2866_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\] net790 _0767_ _0453_
+ VPWR VGND sg13g2_mux2_1
X_4605_ net668 net719 _0035_ VPWR VGND sg13g2_nor2_1
X_2797_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\] net780 _0751_ _0515_
+ VPWR VGND sg13g2_mux2_1
X_4536_ _2165_ net603 _2136_ VPWR VGND sg13g2_nand2_1
X_4467_ _2101_ _0653_ _2088_ VPWR VGND sg13g2_xnor2_1
Xfanout802 net805 net802 VPWR VGND sg13g2_buf_8
X_3418_ VGND VPWR _1069_ _1071_ _1087_ _1085_ sg13g2_a21oi_1
X_4398_ _2043_ _2042_ _0910_ VPWR VGND sg13g2_nand2b_1
X_3349_ videogen.fancy_shader.video_y\[1\] _1030_ _1032_ VPWR VGND sg13g2_and2_1
X_5019_ net206 VGND VPWR _0447_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\]
+ _0104_ sg13g2_dfrbpq_1
XFILLER_27_977 VPWR VGND sg13g2_decap_8
XFILLER_42_11 VPWR VGND sg13g2_fill_2
XFILLER_41_446 VPWR VGND sg13g2_decap_4
XFILLER_9_119 VPWR VGND sg13g2_fill_2
XFILLER_13_159 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_fill_2
XFILLER_21_170 VPWR VGND sg13g2_decap_4
XFILLER_5_303 VPWR VGND sg13g2_fill_2
XFILLER_10_888 VPWR VGND sg13g2_decap_8
XFILLER_3_38 VPWR VGND sg13g2_decap_4
XFILLER_49_513 VPWR VGND sg13g2_decap_8
XFILLER_1_564 VPWR VGND sg13g2_decap_8
XFILLER_18_933 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk_regs clknet_0_clk_regs clknet_3_1__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_17_432 VPWR VGND sg13g2_decap_4
XFILLER_33_903 VPWR VGND sg13g2_decap_8
X_4998__247 VPWR VGND net247 sg13g2_tiehi
X_5024__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_34_1013 VPWR VGND sg13g2_decap_8
X_2720_ net772 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\] _0731_ _0572_
+ VPWR VGND sg13g2_mux2_1
X_2651_ _0685_ _0703_ _0704_ VPWR VGND sg13g2_and2_1
X_2582_ VPWR _0638_ videogen.fancy_shader.video_y\[8\] VGND sg13g2_inv_1
XFILLER_5_881 VPWR VGND sg13g2_decap_8
X_4321_ _1693_ _1974_ net797 _1979_ VPWR VGND sg13g2_nand3_1
X_4252_ VPWR _1914_ _1913_ VGND sg13g2_inv_1
X_3203_ net797 VPWR _0925_ VGND videogen.fancy_shader.video_x\[3\] _0811_ sg13g2_o21ai_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_4183_ _1835_ VPWR _1845_ VGND _1843_ _1844_ sg13g2_o21ai_1
X_3134_ _0863_ tmds_green.n126 _0864_ VPWR VGND sg13g2_xor2_1
XFILLER_27_207 VPWR VGND sg13g2_fill_2
X_3065_ VGND VPWR _0835_ _0847_ net18 _0836_ sg13g2_a21oi_1
X_4981__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_24_969 VPWR VGND sg13g2_decap_8
X_3967_ _1631_ _1632_ _1633_ _1634_ _1635_ VPWR VGND sg13g2_nor4_1
X_2918_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\] _0782_ _0416_
+ VPWR VGND sg13g2_mux2_1
X_3898_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\] net569 _1567_ VPWR
+ VGND sg13g2_nor2_1
X_2849_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\] net780 _0763_ _0466_
+ VPWR VGND sg13g2_mux2_1
X_4953__331 VPWR VGND net331 sg13g2_tiehi
XFILLER_3_829 VPWR VGND sg13g2_decap_8
X_4519_ _2149_ _2134_ _2146_ VPWR VGND sg13g2_xnor2_1
Xfanout632 net640 net632 VPWR VGND sg13g2_buf_8
Xfanout610 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] net610 VPWR VGND
+ sg13g2_buf_8
Xfanout621 net622 net621 VPWR VGND sg13g2_buf_8
Xfanout665 net666 net665 VPWR VGND sg13g2_buf_8
Xfanout643 net646 net643 VPWR VGND sg13g2_buf_8
X_5047__130 VPWR VGND net130 sg13g2_tiehi
Xfanout654 net672 net654 VPWR VGND sg13g2_buf_1
Xfanout676 net682 net676 VPWR VGND sg13g2_buf_1
Xfanout698 net699 net698 VPWR VGND sg13g2_buf_1
Xfanout687 net693 net687 VPWR VGND sg13g2_buf_8
XFILLER_46_549 VPWR VGND sg13g2_decap_8
XFILLER_18_218 VPWR VGND sg13g2_decap_8
XFILLER_18_229 VPWR VGND sg13g2_fill_2
XFILLER_27_730 VPWR VGND sg13g2_decap_8
XFILLER_26_240 VPWR VGND sg13g2_decap_4
X_4960__324 VPWR VGND net324 sg13g2_tiehi
XFILLER_14_413 VPWR VGND sg13g2_fill_2
XFILLER_15_947 VPWR VGND sg13g2_decap_8
XFILLER_41_243 VPWR VGND sg13g2_decap_8
XFILLER_30_917 VPWR VGND sg13g2_decap_8
XFILLER_5_122 VPWR VGND sg13g2_decap_8
XFILLER_45_9 VPWR VGND sg13g2_fill_1
XFILLER_2_873 VPWR VGND sg13g2_decap_8
X_5065__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_49_376 VPWR VGND sg13g2_decap_8
XFILLER_37_527 VPWR VGND sg13g2_fill_2
XFILLER_18_741 VPWR VGND sg13g2_decap_8
XFILLER_33_711 VPWR VGND sg13g2_decap_4
X_4870_ net99 VGND VPWR _0298_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[3\]
+ _0029_ sg13g2_dfrbpq_1
XFILLER_32_221 VPWR VGND sg13g2_fill_1
X_3821_ net616 _1484_ _1489_ _1490_ VPWR VGND sg13g2_nor3_1
XFILLER_32_265 VPWR VGND sg13g2_fill_1
XFILLER_14_980 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_8
X_3752_ net596 _1415_ _1420_ _1421_ VPWR VGND sg13g2_nor3_1
X_3683_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\] net575 _1352_ VPWR
+ VGND sg13g2_nor2_1
X_2703_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\] net760 _0727_ _0585_
+ VPWR VGND sg13g2_mux2_1
X_4937__348 VPWR VGND net348 sg13g2_tiehi
X_2634_ VGND VPWR _0687_ net628 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\]
+ sg13g2_or2_1
X_4304_ _1236_ VPWR _1966_ VGND _1957_ _1958_ sg13g2_o21ai_1
X_4235_ _1881_ _1889_ _1897_ VPWR VGND sg13g2_nor2_1
X_4166_ _1828_ _1009_ _1017_ VPWR VGND sg13g2_xnor2_1
X_3117_ net606 net803 _0852_ VPWR VGND sg13g2_and2_1
X_4097_ _1760_ _1761_ _1762_ VPWR VGND sg13g2_and2_1
X_3048_ _0677_ _0833_ _0835_ VPWR VGND sg13g2_nor2_2
XFILLER_24_711 VPWR VGND sg13g2_fill_1
XFILLER_24_744 VPWR VGND sg13g2_decap_8
XFILLER_36_593 VPWR VGND sg13g2_decap_4
X_4999_ net245 VGND VPWR _0427_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\]
+ _0084_ sg13g2_dfrbpq_1
XFILLER_20_983 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_368 VPWR VGND sg13g2_fill_1
XFILLER_42_530 VPWR VGND sg13g2_fill_1
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_42_552 VPWR VGND sg13g2_decap_8
XFILLER_14_298 VPWR VGND sg13g2_fill_1
XFILLER_31_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_460 VPWR VGND sg13g2_fill_2
XFILLER_11_994 VPWR VGND sg13g2_decap_8
XFILLER_7_976 VPWR VGND sg13g2_decap_8
XFILLER_10_482 VPWR VGND sg13g2_decap_8
X_4020_ net623 _1684_ _1685_ _1687_ _1688_ VPWR VGND sg13g2_nor4_1
X_5147__393 VPWR VGND net393 sg13g2_tiehi
XFILLER_37_313 VPWR VGND sg13g2_fill_2
XFILLER_37_335 VPWR VGND sg13g2_fill_1
X_4943__341 VPWR VGND net341 sg13g2_tiehi
X_4922_ net378 VGND VPWR _0350_ videogen.fancy_shader.n646\[4\] net647 sg13g2_dfrbpq_2
X_4853_ net133 VGND VPWR _0281_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\]
+ _0012_ sg13g2_dfrbpq_1
X_3804_ net623 _1469_ _1470_ _1472_ _1473_ VPWR VGND sg13g2_nor4_1
XFILLER_20_235 VPWR VGND sg13g2_fill_2
X_4784_ net657 net709 _0214_ VPWR VGND sg13g2_nor2_1
X_3735_ _1400_ _1401_ _1402_ _1403_ _1404_ VPWR VGND sg13g2_nor4_1
X_4950__334 VPWR VGND net334 sg13g2_tiehi
Xheichips25_bagel_28 VPWR VGND uio_out[5] sg13g2_tielo
X_3666_ _0646_ _1329_ _1334_ _1335_ VPWR VGND sg13g2_nor3_1
X_2617_ net412 net445 serialize.n433\[1\] VPWR VGND sg13g2_xor2_1
X_3597_ _1076_ _1265_ _1266_ VPWR VGND sg13g2_nor2_1
X_4218_ _1880_ _1806_ _1879_ VPWR VGND sg13g2_xnor2_1
X_5198_ net82 VGND VPWR _0622_ tmds_green.dc_balancing_reg\[4\] net645 sg13g2_dfrbpq_2
X_4149_ _1811_ _1723_ _1809_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_46 VPWR VGND sg13g2_fill_1
XFILLER_18_57 VPWR VGND sg13g2_decap_8
XFILLER_29_858 VPWR VGND sg13g2_decap_8
XFILLER_43_349 VPWR VGND sg13g2_decap_4
XFILLER_36_390 VPWR VGND sg13g2_fill_2
XFILLER_8_707 VPWR VGND sg13g2_decap_8
XFILLER_12_769 VPWR VGND sg13g2_fill_2
Xclkload0 VPWR clkload0/Y clknet_1_1__leaf_clk VGND sg13g2_inv_1
XFILLER_4_946 VPWR VGND sg13g2_decap_8
XFILLER_35_828 VPWR VGND sg13g2_decap_4
XFILLER_34_338 VPWR VGND sg13g2_decap_8
XFILLER_34_349 VPWR VGND sg13g2_fill_1
XFILLER_30_511 VPWR VGND sg13g2_decap_8
XFILLER_30_566 VPWR VGND sg13g2_fill_2
X_3520_ _1189_ _1187_ _1188_ VPWR VGND sg13g2_nand2_1
X_3451_ videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.n646\[6\] _1120_
+ VPWR VGND sg13g2_xor2_1
X_3382_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ _1054_ videogen.test_lut_thingy.gol_counter_reg\[2\] sg13g2_a21oi_1
XFILLER_3_990 VPWR VGND sg13g2_decap_8
X_5121_ net205 VGND VPWR _0545_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\]
+ _0193_ sg13g2_dfrbpq_1
X_5052_ net110 VGND VPWR _0480_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\]
+ _0137_ sg13g2_dfrbpq_1
XFILLER_38_633 VPWR VGND sg13g2_decap_8
X_4003_ _1670_ VPWR _1671_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\]
+ net579 sg13g2_o21ai_1
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_26_839 VPWR VGND sg13g2_decap_8
X_4905_ net40 VGND VPWR _0333_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\]
+ net630 sg13g2_dfrbpq_1
XFILLER_21_511 VPWR VGND sg13g2_fill_1
X_4836_ net156 VGND VPWR _0265_ clockdiv.q1 clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_14_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_599 VPWR VGND sg13g2_fill_1
X_4767_ net667 net720 _0197_ VPWR VGND sg13g2_nor2_1
X_3718_ _1383_ _1384_ _1385_ _1386_ _1387_ VPWR VGND sg13g2_nor4_1
X_4698_ net679 net731 _0128_ VPWR VGND sg13g2_nor2_1
XFILLER_20_58 VPWR VGND sg13g2_fill_1
X_3649_ net617 VPWR _1318_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\]
+ net590 sg13g2_o21ai_1
XFILLER_1_949 VPWR VGND sg13g2_decap_8
Xhold12 serialize.n414\[3\] VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold23 serialize.n417\[0\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold34 serialize.n414\[4\] VPWR VGND net439 sg13g2_dlygate4sd3_1
XFILLER_28_143 VPWR VGND sg13g2_fill_1
XFILLER_45_99 VPWR VGND sg13g2_decap_4
XFILLER_45_66 VPWR VGND sg13g2_decap_8
XFILLER_25_872 VPWR VGND sg13g2_decap_8
XFILLER_31_319 VPWR VGND sg13g2_fill_1
XFILLER_40_831 VPWR VGND sg13g2_decap_4
XFILLER_0_971 VPWR VGND sg13g2_decap_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
XFILLER_35_636 VPWR VGND sg13g2_decap_4
XFILLER_37_1000 VPWR VGND sg13g2_decap_8
XFILLER_16_861 VPWR VGND sg13g2_decap_8
X_4940__344 VPWR VGND net344 sg13g2_tiehi
XFILLER_15_360 VPWR VGND sg13g2_decap_4
XFILLER_22_308 VPWR VGND sg13g2_fill_2
X_2951_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\] _0791_ _0392_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_853 VPWR VGND sg13g2_fill_1
X_2882_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\] net753 _0774_ _0444_
+ VPWR VGND sg13g2_mux2_1
X_4621_ net662 net714 _0051_ VPWR VGND sg13g2_nor2_1
X_4552_ _2180_ _2176_ _2181_ VPWR VGND sg13g2_xor2_1
X_4483_ _0856_ _2111_ _2116_ _2117_ VPWR VGND sg13g2_nor3_1
X_3503_ _1148_ _1169_ _1171_ _1172_ VPWR VGND sg13g2_or3_1
X_5034__176 VPWR VGND net176 sg13g2_tiehi
X_3434_ VGND VPWR _1102_ _1103_ videogen.fancy_shader.n646\[7\] videogen.fancy_shader.video_y\[7\]
+ sg13g2_a21oi_2
X_4878__90 VPWR VGND net90 sg13g2_tiehi
X_3365_ net745 _1042_ _1044_ _0360_ VPWR VGND sg13g2_nor3_1
X_5104_ net275 VGND VPWR _0528_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\]
+ _0176_ sg13g2_dfrbpq_1
X_3296_ _0988_ net608 videogen.fancy_shader.n646\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_39_964 VPWR VGND sg13g2_fill_1
X_5035_ net174 VGND VPWR _0463_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\]
+ _0120_ sg13g2_dfrbpq_1
XFILLER_39_997 VPWR VGND sg13g2_decap_8
XFILLER_38_496 VPWR VGND sg13g2_decap_4
XFILLER_41_628 VPWR VGND sg13g2_fill_2
XFILLER_13_308 VPWR VGND sg13g2_fill_1
XFILLER_21_330 VPWR VGND sg13g2_fill_2
XFILLER_22_831 VPWR VGND sg13g2_fill_2
XFILLER_22_897 VPWR VGND sg13g2_decap_8
XFILLER_31_24 VPWR VGND sg13g2_fill_2
X_4819_ net688 net740 _0249_ VPWR VGND sg13g2_nor2_1
Xoutput13 net13 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_724 VPWR VGND sg13g2_decap_8
XFILLER_0_234 VPWR VGND sg13g2_fill_1
XFILLER_0_267 VPWR VGND sg13g2_fill_1
Xclkbuf_3_0__f_clk_regs clknet_0_clk_regs clknet_3_0__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_4846__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_44_444 VPWR VGND sg13g2_decap_4
XFILLER_16_146 VPWR VGND sg13g2_fill_2
XFILLER_16_168 VPWR VGND sg13g2_fill_2
XFILLER_32_639 VPWR VGND sg13g2_decap_8
XFILLER_25_691 VPWR VGND sg13g2_fill_1
XFILLER_31_138 VPWR VGND sg13g2_decap_8
XFILLER_12_341 VPWR VGND sg13g2_decap_4
XFILLER_12_352 VPWR VGND sg13g2_decap_8
XFILLER_8_334 VPWR VGND sg13g2_fill_2
XFILLER_9_846 VPWR VGND sg13g2_fill_2
XFILLER_9_868 VPWR VGND sg13g2_decap_8
XFILLER_12_374 VPWR VGND sg13g2_decap_8
X_3150_ _0879_ _0663_ _0875_ VPWR VGND sg13g2_nand2_1
X_3081_ net428 blue_tmds_par\[0\] net697 serialize.n429\[0\] VPWR VGND sg13g2_mux2_1
XFILLER_39_227 VPWR VGND sg13g2_fill_1
X_4875__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_35_444 VPWR VGND sg13g2_decap_4
XFILLER_35_466 VPWR VGND sg13g2_fill_2
XFILLER_22_105 VPWR VGND sg13g2_decap_4
X_3983_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\] net580 _1651_ VPWR
+ VGND sg13g2_nor2_1
X_2934_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\] net762 _0785_ _0403_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_672 VPWR VGND sg13g2_fill_1
X_2865_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\] net779 _0767_ _0454_
+ VPWR VGND sg13g2_mux2_1
X_4604_ net683 net734 _0034_ VPWR VGND sg13g2_nor2_1
X_2796_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\] net768 _0751_ _0516_
+ VPWR VGND sg13g2_mux2_1
X_4535_ _2164_ tmds_blue.dc_balancing_reg\[3\] _2140_ VPWR VGND sg13g2_xnor2_1
X_5186__227 VPWR VGND net227 sg13g2_tiehi
X_4466_ net571 _2100_ _0620_ VPWR VGND sg13g2_nor2_1
X_4916__390 VPWR VGND net390 sg13g2_tiehi
Xfanout803 net804 net803 VPWR VGND sg13g2_buf_8
X_3417_ _1086_ _1069_ _1071_ _1085_ VPWR VGND sg13g2_and3_1
X_4397_ _2042_ _2019_ _2035_ VPWR VGND sg13g2_xnor2_1
X_3348_ _1030_ _1031_ _0356_ VPWR VGND sg13g2_nor2_1
X_5086__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_39_761 VPWR VGND sg13g2_fill_2
XFILLER_39_750 VPWR VGND sg13g2_decap_8
X_3279_ _0818_ _0975_ _0976_ _0334_ VPWR VGND sg13g2_nor3_1
XFILLER_27_901 VPWR VGND sg13g2_fill_2
X_5018_ net208 VGND VPWR _0446_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\]
+ _0103_ sg13g2_dfrbpq_1
XFILLER_38_271 VPWR VGND sg13g2_decap_8
XFILLER_26_13 VPWR VGND sg13g2_fill_1
XFILLER_26_24 VPWR VGND sg13g2_fill_2
XFILLER_27_956 VPWR VGND sg13g2_decap_8
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_13_149 VPWR VGND sg13g2_decap_4
XFILLER_10_834 VPWR VGND sg13g2_fill_1
XFILLER_10_845 VPWR VGND sg13g2_fill_1
XFILLER_6_805 VPWR VGND sg13g2_fill_1
XFILLER_1_543 VPWR VGND sg13g2_decap_8
X_5128__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_49_569 VPWR VGND sg13g2_decap_8
XFILLER_18_912 VPWR VGND sg13g2_decap_8
XFILLER_17_400 VPWR VGND sg13g2_fill_1
X_4872__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_44_274 VPWR VGND sg13g2_fill_1
XFILLER_18_989 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_9_610 VPWR VGND sg13g2_fill_1
XFILLER_20_609 VPWR VGND sg13g2_fill_2
XFILLER_13_672 VPWR VGND sg13g2_fill_1
XFILLER_8_142 VPWR VGND sg13g2_fill_2
XFILLER_12_182 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_fill_1
X_2650_ net593 net583 _0703_ VPWR VGND sg13g2_nor2_1
X_2581_ VPWR _0637_ videogen.fancy_shader.video_y\[9\] VGND sg13g2_inv_1
X_4320_ VGND VPWR _1972_ _1978_ _0382_ net747 sg13g2_a21oi_1
X_4251_ _1910_ _1902_ _1913_ VPWR VGND sg13g2_xor2_1
X_3202_ net750 _0811_ _0924_ _0301_ VPWR VGND sg13g2_nor3_1
XFILLER_41_1007 VPWR VGND sg13g2_decap_8
X_4182_ VGND VPWR _1820_ _1833_ _1844_ _1834_ sg13g2_a21oi_1
X_3133_ _0862_ VPWR _0863_ VGND _0855_ _0859_ sg13g2_o21ai_1
X_3064_ _0843_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0847_ VPWR VGND
+ sg13g2_xor2_1
XFILLER_36_786 VPWR VGND sg13g2_decap_8
X_5003__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_24_948 VPWR VGND sg13g2_decap_8
X_3966_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\] net584 _1634_ VPWR
+ VGND sg13g2_nor2_1
X_2917_ _0782_ _0720_ _0781_ VPWR VGND sg13g2_nand2_2
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_3897_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\] net591 _1566_ VPWR
+ VGND sg13g2_nor2_1
X_2848_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\] net768 _0763_ _0467_
+ VPWR VGND sg13g2_mux2_1
XFILLER_3_808 VPWR VGND sg13g2_decap_8
X_2779_ _0712_ _0745_ _0748_ VPWR VGND sg13g2_nor2_2
X_4518_ _2148_ net602 _2147_ VPWR VGND sg13g2_nand2_1
XFILLER_2_329 VPWR VGND sg13g2_decap_8
X_4449_ net600 net599 tmds_green.n126 _2084_ VPWR VGND sg13g2_nor3_1
Xfanout600 net601 net600 VPWR VGND sg13g2_buf_8
Xfanout611 net613 net611 VPWR VGND sg13g2_buf_8
Xfanout633 net640 net633 VPWR VGND sg13g2_buf_8
Xfanout622 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\] net622 VPWR VGND
+ sg13g2_buf_8
Xfanout666 net672 net666 VPWR VGND sg13g2_buf_8
Xfanout655 net656 net655 VPWR VGND sg13g2_buf_8
Xfanout644 net646 net644 VPWR VGND sg13g2_buf_8
Xfanout699 net700 net699 VPWR VGND sg13g2_buf_8
Xfanout688 net692 net688 VPWR VGND sg13g2_buf_8
XFILLER_37_12 VPWR VGND sg13g2_decap_4
Xfanout677 net682 net677 VPWR VGND sg13g2_buf_8
XFILLER_37_89 VPWR VGND sg13g2_fill_1
X_4843__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_15_926 VPWR VGND sg13g2_decap_8
XFILLER_41_233 VPWR VGND sg13g2_fill_2
XFILLER_14_425 VPWR VGND sg13g2_decap_4
XFILLER_42_767 VPWR VGND sg13g2_fill_1
XFILLER_41_266 VPWR VGND sg13g2_decap_8
X_5054__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_10_642 VPWR VGND sg13g2_decap_4
XFILLER_10_675 VPWR VGND sg13g2_decap_4
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_2_852 VPWR VGND sg13g2_decap_8
X_4850__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_38_9 VPWR VGND sg13g2_fill_1
X_3820_ net623 _1485_ _1487_ _1488_ _1489_ VPWR VGND sg13g2_nor4_1
XFILLER_21_929 VPWR VGND sg13g2_decap_8
XFILLER_20_439 VPWR VGND sg13g2_fill_2
X_3751_ net622 _1416_ _1417_ _1419_ _1420_ VPWR VGND sg13g2_nor4_1
X_2702_ _0719_ _0726_ _0727_ VPWR VGND sg13g2_nor2_2
X_3682_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\] net586 _1351_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_484 VPWR VGND sg13g2_decap_8
XFILLER_9_495 VPWR VGND sg13g2_fill_1
X_2633_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\] net628 _0686_ VPWR VGND
+ sg13g2_nor2_1
X_4303_ _1865_ _1235_ _1964_ _1965_ VPWR VGND sg13g2_a21o_1
X_4234_ _1893_ _1895_ _1892_ _1896_ VPWR VGND sg13g2_nand3_1
X_4165_ _1827_ _1821_ _1826_ VPWR VGND sg13g2_xnor2_1
X_3116_ _0822_ _0825_ _0000_ VPWR VGND sg13g2_nor2_1
XFILLER_28_517 VPWR VGND sg13g2_fill_2
X_4096_ _1739_ VPWR _1761_ VGND _1744_ _1759_ sg13g2_o21ai_1
X_3047_ _0829_ _0831_ _0834_ VPWR VGND sg13g2_nor2_1
XFILLER_24_701 VPWR VGND sg13g2_fill_2
X_4998_ net247 VGND VPWR _0426_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\]
+ _0083_ sg13g2_dfrbpq_1
XFILLER_23_36 VPWR VGND sg13g2_decap_4
XFILLER_20_962 VPWR VGND sg13g2_decap_8
X_3949_ net622 _1613_ _1615_ _1616_ _1617_ VPWR VGND sg13g2_nor4_1
X_5207__403 VPWR VGND net403 sg13g2_tiehi
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_15_789 VPWR VGND sg13g2_fill_2
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_955 VPWR VGND sg13g2_decap_8
XFILLER_49_185 VPWR VGND sg13g2_decap_8
XFILLER_37_347 VPWR VGND sg13g2_fill_2
XFILLER_46_881 VPWR VGND sg13g2_decap_8
X_4921_ net380 VGND VPWR _0349_ videogen.fancy_shader.n646\[3\] net647 sg13g2_dfrbpq_2
XFILLER_18_583 VPWR VGND sg13g2_decap_8
XFILLER_33_531 VPWR VGND sg13g2_decap_8
XFILLER_45_391 VPWR VGND sg13g2_decap_8
X_4852_ net135 VGND VPWR _0280_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\]
+ _0011_ sg13g2_dfrbpq_1
XFILLER_33_564 VPWR VGND sg13g2_decap_8
X_3803_ _1471_ VPWR _1472_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\]
+ net589 sg13g2_o21ai_1
XFILLER_21_737 VPWR VGND sg13g2_decap_8
X_4783_ net658 net710 _0213_ VPWR VGND sg13g2_nor2_1
XFILLER_21_748 VPWR VGND sg13g2_fill_1
X_3734_ net625 VPWR _1403_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\]
+ net569 sg13g2_o21ai_1
X_3665_ _1330_ _1331_ _1332_ _1333_ _1334_ VPWR VGND sg13g2_nor4_1
X_2616_ _0671_ serialize.bit_cnt\[1\] net412 VPWR VGND sg13g2_nand2_1
Xheichips25_bagel_29 VPWR VGND uio_out[6] sg13g2_tielo
X_3596_ VGND VPWR _1250_ _1264_ _1265_ _1261_ sg13g2_a21oi_1
X_4217_ _1154_ _1155_ _1145_ _1879_ VPWR VGND _1876_ sg13g2_nand4_1
X_5197_ net108 VGND VPWR _0621_ tmds_green.dc_balancing_reg\[3\] net645 sg13g2_dfrbpq_1
X_4148_ _1809_ _1723_ _1810_ VPWR VGND sg13g2_xor2_1
XFILLER_43_317 VPWR VGND sg13g2_fill_2
X_4079_ VPWR _1744_ _1743_ VGND sg13g2_inv_1
XFILLER_43_328 VPWR VGND sg13g2_fill_2
XFILLER_24_520 VPWR VGND sg13g2_decap_8
XFILLER_34_13 VPWR VGND sg13g2_decap_4
X_5159__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_12_704 VPWR VGND sg13g2_fill_1
XFILLER_24_531 VPWR VGND sg13g2_fill_1
XFILLER_34_46 VPWR VGND sg13g2_decap_8
XFILLER_34_57 VPWR VGND sg13g2_fill_1
XFILLER_34_79 VPWR VGND sg13g2_fill_1
XFILLER_11_236 VPWR VGND sg13g2_decap_8
Xclkload1 VPWR clkload1/Y clknet_3_1__leaf_clk_regs VGND sg13g2_inv_1
XFILLER_20_770 VPWR VGND sg13g2_decap_8
XFILLER_4_925 VPWR VGND sg13g2_decap_8
XFILLER_3_468 VPWR VGND sg13g2_decap_8
XFILLER_42_361 VPWR VGND sg13g2_fill_2
X_3450_ _1119_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.video_x\[6\]
+ VPWR VGND sg13g2_nand2_1
X_3381_ VGND VPWR videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ _0367_ _1053_ sg13g2_a21oi_1
X_5120_ net209 VGND VPWR _0544_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\]
+ _0192_ sg13g2_dfrbpq_1
X_5051_ net114 VGND VPWR _0479_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\]
+ _0136_ sg13g2_dfrbpq_1
X_4002_ VGND VPWR _1670_ net566 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\]
+ sg13g2_or2_1
XFILLER_37_122 VPWR VGND sg13g2_decap_4
XFILLER_26_818 VPWR VGND sg13g2_decap_8
X_4904_ net42 VGND VPWR _0332_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\]
+ net630 sg13g2_dfrbpq_1
XFILLER_21_556 VPWR VGND sg13g2_decap_8
X_4835_ net158 VGND VPWR _0264_ tmds_blue.dc_balancing_reg\[0\] net643 sg13g2_dfrbpq_1
XFILLER_14_1001 VPWR VGND sg13g2_decap_8
XFILLER_21_567 VPWR VGND sg13g2_fill_1
X_4766_ net667 net720 _0196_ VPWR VGND sg13g2_nor2_1
X_3717_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\] net557 _1386_ VPWR
+ VGND sg13g2_nor2_1
X_5189__203 VPWR VGND net203 sg13g2_tiehi
X_4697_ net679 net731 _0127_ VPWR VGND sg13g2_nor2_1
X_3648_ _1313_ _1314_ _1315_ _1316_ _1317_ VPWR VGND sg13g2_nor4_1
X_3579_ _1146_ _1247_ _1248_ VPWR VGND sg13g2_and2_1
XFILLER_1_928 VPWR VGND sg13g2_decap_8
XFILLER_48_409 VPWR VGND sg13g2_decap_8
Xhold13 serialize.n414\[5\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold35 serialize.n417\[1\] VPWR VGND net440 sg13g2_dlygate4sd3_1
Xhold24 serialize.n414\[6\] VPWR VGND net429 sg13g2_dlygate4sd3_1
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_122 VPWR VGND sg13g2_fill_1
XFILLER_29_634 VPWR VGND sg13g2_fill_1
XFILLER_17_829 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_4
XFILLER_45_34 VPWR VGND sg13g2_fill_1
X_4926__370 VPWR VGND net370 sg13g2_tiehi
XFILLER_25_851 VPWR VGND sg13g2_decap_8
XFILLER_40_887 VPWR VGND sg13g2_fill_2
XFILLER_8_527 VPWR VGND sg13g2_decap_8
XFILLER_12_589 VPWR VGND sg13g2_decap_8
XFILLER_4_700 VPWR VGND sg13g2_fill_2
XFILLER_4_744 VPWR VGND sg13g2_fill_1
XFILLER_3_221 VPWR VGND sg13g2_fill_1
XFILLER_0_950 VPWR VGND sg13g2_decap_8
XFILLER_48_921 VPWR VGND sg13g2_decap_8
XFILLER_13_8 VPWR VGND sg13g2_fill_2
XFILLER_48_998 VPWR VGND sg13g2_decap_8
XFILLER_47_453 VPWR VGND sg13g2_decap_4
XFILLER_34_136 VPWR VGND sg13g2_fill_2
XFILLER_43_670 VPWR VGND sg13g2_fill_2
X_5071__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_15_350 VPWR VGND sg13g2_decap_4
X_2950_ _0791_ _0781_ VPWR VGND _0707_ sg13g2_nand2b_2
X_2881_ _0714_ _0726_ _0774_ VPWR VGND sg13g2_nor2_2
X_4620_ net661 net713 _0050_ VPWR VGND sg13g2_nor2_1
X_4551_ _2178_ _2164_ _2180_ VPWR VGND sg13g2_xor2_1
X_4482_ _0863_ _2115_ _2116_ VPWR VGND sg13g2_nor2_1
X_3502_ _1171_ _1090_ _1158_ VPWR VGND sg13g2_nand2_1
X_4834__261 VPWR VGND net261 sg13g2_tiehi
X_3433_ VGND VPWR _0639_ _0642_ _1102_ _1098_ sg13g2_a21oi_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
X_5103_ net279 VGND VPWR _0527_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\]
+ _0175_ sg13g2_dfrbpq_1
X_3364_ videogen.fancy_shader.video_y\[4\] _1041_ _1044_ VPWR VGND sg13g2_and2_1
XFILLER_32_0 VPWR VGND sg13g2_decap_8
X_3295_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_y\[1\] _0987_
+ VPWR VGND sg13g2_xor2_1
XFILLER_39_932 VPWR VGND sg13g2_decap_8
X_5034_ net176 VGND VPWR _0462_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\]
+ _0119_ sg13g2_dfrbpq_1
XFILLER_39_976 VPWR VGND sg13g2_decap_8
XFILLER_41_607 VPWR VGND sg13g2_decap_8
XFILLER_25_158 VPWR VGND sg13g2_fill_2
XFILLER_34_670 VPWR VGND sg13g2_fill_2
X_4818_ net688 net735 _0248_ VPWR VGND sg13g2_nor2_1
X_4991__265 VPWR VGND net265 sg13g2_tiehi
X_4749_ net673 net725 _0179_ VPWR VGND sg13g2_nor2_1
Xoutput14 net14 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_0_246 VPWR VGND sg13g2_decap_8
XFILLER_0_213 VPWR VGND sg13g2_decap_8
XFILLER_1_747 VPWR VGND sg13g2_fill_1
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_29_431 VPWR VGND sg13g2_decap_8
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_17_626 VPWR VGND sg13g2_decap_8
XFILLER_16_125 VPWR VGND sg13g2_decap_8
XFILLER_32_618 VPWR VGND sg13g2_decap_8
XFILLER_9_803 VPWR VGND sg13g2_fill_1
XFILLER_8_313 VPWR VGND sg13g2_fill_1
XFILLER_13_898 VPWR VGND sg13g2_decap_8
X_4970__305 VPWR VGND net305 sg13g2_tiehi
XFILLER_4_574 VPWR VGND sg13g2_decap_8
X_3080_ VGND VPWR serialize.n431\[6\] net700 net419 sg13g2_or2_1
XFILLER_36_924 VPWR VGND sg13g2_fill_1
XFILLER_35_412 VPWR VGND sg13g2_fill_1
X_3982_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\] net590 _1650_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_16_681 VPWR VGND sg13g2_fill_1
X_2933_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\] net753 _0785_ _0404_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_651 VPWR VGND sg13g2_fill_2
X_2864_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\] net767 _0767_ _0455_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_684 VPWR VGND sg13g2_decap_4
X_2795_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\] net758 _0751_ _0517_
+ VPWR VGND sg13g2_mux2_1
X_4603_ net660 net712 _0033_ VPWR VGND sg13g2_nor2_1
XFILLER_30_183 VPWR VGND sg13g2_decap_4
X_4534_ _2160_ _2163_ _0625_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_891 VPWR VGND sg13g2_decap_8
XFILLER_7_82 VPWR VGND sg13g2_decap_8
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
X_4465_ _2100_ _0860_ _2099_ VPWR VGND sg13g2_xnor2_1
Xfanout804 net805 net804 VPWR VGND sg13g2_buf_8
X_3416_ _1085_ _1084_ _1083_ VPWR VGND sg13g2_nand2b_1
X_4396_ VPWR _2041_ _2040_ VGND sg13g2_inv_1
X_3347_ net797 VPWR _1031_ VGND net608 _0922_ sg13g2_o21ai_1
X_5017_ net210 VGND VPWR _0445_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\]
+ _0102_ sg13g2_dfrbpq_1
X_3278_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0807_ _0976_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_39_784 VPWR VGND sg13g2_fill_1
XFILLER_38_250 VPWR VGND sg13g2_decap_8
XFILLER_27_935 VPWR VGND sg13g2_decap_8
XFILLER_26_36 VPWR VGND sg13g2_decap_8
XFILLER_41_415 VPWR VGND sg13g2_decap_4
XFILLER_14_629 VPWR VGND sg13g2_fill_2
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_42_46 VPWR VGND sg13g2_decap_4
XFILLER_21_150 VPWR VGND sg13g2_fill_2
XFILLER_22_695 VPWR VGND sg13g2_decap_8
XFILLER_42_79 VPWR VGND sg13g2_fill_1
XFILLER_5_338 VPWR VGND sg13g2_fill_2
XFILLER_3_18 VPWR VGND sg13g2_fill_1
XFILLER_1_522 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_decap_8
XFILLER_29_261 VPWR VGND sg13g2_fill_2
XFILLER_44_231 VPWR VGND sg13g2_fill_2
XFILLER_18_968 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
X_5098__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_41_993 VPWR VGND sg13g2_decap_8
XFILLER_9_644 VPWR VGND sg13g2_decap_8
XFILLER_13_684 VPWR VGND sg13g2_decap_4
XFILLER_9_666 VPWR VGND sg13g2_decap_4
XFILLER_9_699 VPWR VGND sg13g2_fill_1
X_2580_ VPWR _0636_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[0\] VGND
+ sg13g2_inv_1
X_4250_ VGND VPWR _1904_ _1907_ _1912_ _1911_ sg13g2_a21oi_1
X_3201_ videogen.fancy_shader.video_x\[2\] _0810_ _0924_ VPWR VGND sg13g2_nor2_1
X_4181_ VPWR _1843_ _1842_ VGND sg13g2_inv_1
X_3132_ _0862_ tmds_green.dc_balancing_reg\[4\] net601 VPWR VGND sg13g2_nand2b_1
X_3063_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\]
+ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0846_ VPWR VGND _0840_ sg13g2_nand4_1
XFILLER_27_209 VPWR VGND sg13g2_fill_1
XFILLER_24_927 VPWR VGND sg13g2_decap_8
X_3965_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\] net551 _1633_ VPWR
+ VGND sg13g2_nor2_1
X_3896_ net612 _1553_ _1564_ _1565_ VPWR VGND sg13g2_nor3_1
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_2916_ net546 _0770_ _0781_ VPWR VGND sg13g2_and2_1
X_2847_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\] net758 _0763_ _0468_
+ VPWR VGND sg13g2_mux2_1
X_2778_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\] _0747_ _0530_
+ VPWR VGND sg13g2_mux2_1
X_4517_ _2134_ _2146_ _2147_ VPWR VGND sg13g2_nor2_1
X_4448_ net599 tmds_green.n126 _2083_ VPWR VGND sg13g2_nor2_1
Xfanout601 tmds_green.n100 net601 VPWR VGND sg13g2_buf_2
Xfanout612 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] net612 VPWR VGND
+ sg13g2_buf_8
Xfanout623 net627 net623 VPWR VGND sg13g2_buf_8
Xfanout645 net646 net645 VPWR VGND sg13g2_buf_1
Xfanout634 net640 net634 VPWR VGND sg13g2_buf_8
Xfanout656 net659 net656 VPWR VGND sg13g2_buf_8
X_4379_ _2024_ _0666_ _2023_ VPWR VGND sg13g2_xnor2_1
Xfanout667 net671 net667 VPWR VGND sg13g2_buf_8
Xfanout689 net692 net689 VPWR VGND sg13g2_buf_2
Xfanout678 net682 net678 VPWR VGND sg13g2_buf_1
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_fill_1
XFILLER_39_592 VPWR VGND sg13g2_fill_2
XFILLER_15_905 VPWR VGND sg13g2_decap_8
XFILLER_27_765 VPWR VGND sg13g2_fill_2
X_4909__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_10_610 VPWR VGND sg13g2_fill_2
XFILLER_23_993 VPWR VGND sg13g2_decap_8
XFILLER_6_625 VPWR VGND sg13g2_decap_4
XFILLER_6_658 VPWR VGND sg13g2_decap_4
XFILLER_2_831 VPWR VGND sg13g2_decap_8
XFILLER_49_345 VPWR VGND sg13g2_decap_8
XFILLER_49_334 VPWR VGND sg13g2_fill_1
XFILLER_49_367 VPWR VGND sg13g2_decap_4
XFILLER_37_529 VPWR VGND sg13g2_fill_1
XFILLER_45_551 VPWR VGND sg13g2_decap_8
XFILLER_17_264 VPWR VGND sg13g2_fill_2
XFILLER_18_765 VPWR VGND sg13g2_fill_2
XFILLER_27_90 VPWR VGND sg13g2_decap_4
XFILLER_32_212 VPWR VGND sg13g2_decap_8
XFILLER_21_908 VPWR VGND sg13g2_decap_8
XFILLER_32_256 VPWR VGND sg13g2_fill_2
XFILLER_20_418 VPWR VGND sg13g2_fill_1
X_3750_ _1418_ VPWR _1419_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\]
+ net555 sg13g2_o21ai_1
XFILLER_32_289 VPWR VGND sg13g2_decap_4
XFILLER_9_441 VPWR VGND sg13g2_decap_4
XFILLER_13_492 VPWR VGND sg13g2_fill_2
X_2701_ _0704_ _0706_ net619 _0726_ VPWR VGND sg13g2_nand3_1
X_3681_ net615 VPWR _1350_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\]
+ net563 sg13g2_o21ai_1
X_2632_ _0685_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] _0684_ VPWR VGND
+ sg13g2_nand2_2
X_4302_ _1860_ _1864_ _1964_ VPWR VGND sg13g2_and2_1
X_4233_ _1877_ _1888_ _1895_ VPWR VGND sg13g2_nor2b_1
X_4164_ VGND VPWR _1817_ _1825_ _1826_ _1822_ sg13g2_a21oi_1
X_3115_ _0823_ _0851_ _0001_ VPWR VGND sg13g2_nor2_1
X_4095_ _1739_ _1744_ _1759_ _1760_ VPWR VGND sg13g2_or3_1
X_3046_ _0829_ _0830_ _0831_ _0832_ _0833_ VPWR VGND sg13g2_nor4_1
XFILLER_36_562 VPWR VGND sg13g2_fill_1
XFILLER_23_212 VPWR VGND sg13g2_fill_2
XFILLER_12_919 VPWR VGND sg13g2_decap_8
X_4997_ net249 VGND VPWR _0425_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\]
+ _0082_ sg13g2_dfrbpq_1
XFILLER_17_1010 VPWR VGND sg13g2_decap_8
XFILLER_20_941 VPWR VGND sg13g2_decap_8
X_3948_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\] net555 _1616_ VPWR
+ VGND sg13g2_nor2_1
X_3879_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\] net563 _1548_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_2_138 VPWR VGND sg13g2_fill_1
XFILLER_2_149 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_24_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_827 VPWR VGND sg13g2_fill_1
XFILLER_19_507 VPWR VGND sg13g2_decap_4
XFILLER_46_337 VPWR VGND sg13g2_decap_4
XFILLER_27_540 VPWR VGND sg13g2_decap_8
XFILLER_42_521 VPWR VGND sg13g2_decap_4
XFILLER_14_245 VPWR VGND sg13g2_decap_4
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_7_934 VPWR VGND sg13g2_decap_8
X_4936__350 VPWR VGND net350 sg13g2_tiehi
XFILLER_2_650 VPWR VGND sg13g2_fill_1
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_164 VPWR VGND sg13g2_decap_8
XFILLER_37_326 VPWR VGND sg13g2_decap_8
XFILLER_46_860 VPWR VGND sg13g2_decap_8
X_4920_ net382 VGND VPWR _0348_ videogen.fancy_shader.n646\[2\] net647 sg13g2_dfrbpq_2
X_4851_ net137 VGND VPWR _0279_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\]
+ _0010_ sg13g2_dfrbpq_1
X_3802_ VGND VPWR _1471_ net566 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\]
+ sg13g2_or2_1
XFILLER_33_576 VPWR VGND sg13g2_fill_1
XFILLER_20_237 VPWR VGND sg13g2_fill_1
X_4782_ net675 net727 _0212_ VPWR VGND sg13g2_nor2_1
X_3733_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\] net559 _1402_ VPWR
+ VGND sg13g2_nor2_1
X_3664_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\] net573 _1333_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_282 VPWR VGND sg13g2_decap_8
X_2615_ VPWR _0670_ net418 VGND sg13g2_inv_1
Xheichips25_bagel_19 VPWR VGND uio_oe[0] sg13g2_tielo
X_3595_ _1076_ _1259_ _1262_ _1264_ VPWR VGND sg13g2_nor3_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
XFILLER_0_609 VPWR VGND sg13g2_decap_8
X_5196_ net124 VGND VPWR _0620_ tmds_green.dc_balancing_reg\[2\] net645 sg13g2_dfrbpq_1
X_4216_ _1878_ _1145_ _1876_ VPWR VGND sg13g2_nand2_1
X_4147_ _1160_ _1806_ _1809_ VPWR VGND sg13g2_nor2_2
XFILLER_29_838 VPWR VGND sg13g2_fill_1
XFILLER_18_37 VPWR VGND sg13g2_decap_8
XFILLER_43_307 VPWR VGND sg13g2_fill_2
X_4078_ _1743_ _1707_ _1742_ VPWR VGND sg13g2_nand2_1
X_3029_ _0825_ net796 _0824_ VPWR VGND sg13g2_nand2_1
XFILLER_36_370 VPWR VGND sg13g2_decap_8
X_5202__389 VPWR VGND net389 sg13g2_tiehi
XFILLER_34_25 VPWR VGND sg13g2_decap_8
XFILLER_34_36 VPWR VGND sg13g2_fill_2
XFILLER_36_392 VPWR VGND sg13g2_fill_1
Xclkload2 VPWR clkload2/Y clknet_3_3__leaf_clk_regs VGND sg13g2_inv_1
XFILLER_4_904 VPWR VGND sg13g2_decap_8
XFILLER_47_613 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_46_156 VPWR VGND sg13g2_fill_2
XFILLER_46_189 VPWR VGND sg13g2_fill_1
XFILLER_42_340 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_15_587 VPWR VGND sg13g2_fill_1
XFILLER_30_524 VPWR VGND sg13g2_fill_1
XFILLER_30_568 VPWR VGND sg13g2_fill_1
XFILLER_7_775 VPWR VGND sg13g2_fill_2
XFILLER_7_753 VPWR VGND sg13g2_fill_2
X_3380_ net796 VPWR _1053_ VGND videogen.test_lut_thingy.gol_counter_reg\[0\] videogen.test_lut_thingy.gol_counter_reg\[1\]
+ sg13g2_o21ai_1
X_5050_ net118 VGND VPWR _0478_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\]
+ _0135_ sg13g2_dfrbpq_1
X_4001_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\] net557 _1669_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_37_178 VPWR VGND sg13g2_decap_4
X_4903_ net44 VGND VPWR _0331_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\]
+ net630 sg13g2_dfrbpq_1
XFILLER_33_340 VPWR VGND sg13g2_decap_4
X_4834_ net261 VGND VPWR _0263_ tmds_green.dc_balancing_reg\[0\] net645 sg13g2_dfrbpq_1
X_4765_ net662 net714 _0195_ VPWR VGND sg13g2_nor2_1
X_3716_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\] net566 _1385_ VPWR
+ VGND sg13g2_nor2_1
X_4696_ net680 net730 _0126_ VPWR VGND sg13g2_nor2_1
X_3647_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\] net580 _1316_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_1_907 VPWR VGND sg13g2_decap_8
X_3578_ _1139_ _1148_ _1173_ _1247_ VPWR VGND sg13g2_mux2_1
XFILLER_0_428 VPWR VGND sg13g2_decap_8
Xhold14 serialize.n420\[6\] VPWR VGND net419 sg13g2_dlygate4sd3_1
XFILLER_0_439 VPWR VGND sg13g2_decap_8
Xhold36 serialize.n411\[1\] VPWR VGND net441 sg13g2_dlygate4sd3_1
Xhold25 serialize.n411\[6\] VPWR VGND net430 sg13g2_dlygate4sd3_1
X_5248_ net802 VGND VPWR serialize.n427\[9\] serialize.n411\[7\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_69 VPWR VGND sg13g2_fill_2
X_5179_ net381 VGND VPWR _0603_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\]
+ _0251_ sg13g2_dfrbpq_1
XFILLER_21_1006 VPWR VGND sg13g2_decap_8
XFILLER_29_657 VPWR VGND sg13g2_fill_2
XFILLER_16_307 VPWR VGND sg13g2_decap_8
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_12_568 VPWR VGND sg13g2_fill_1
XFILLER_12_579 VPWR VGND sg13g2_decap_4
XFILLER_4_712 VPWR VGND sg13g2_fill_2
XFILLER_3_266 VPWR VGND sg13g2_decap_8
XFILLER_3_288 VPWR VGND sg13g2_decap_4
XFILLER_48_900 VPWR VGND sg13g2_decap_8
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_19_156 VPWR VGND sg13g2_decap_4
XFILLER_35_627 VPWR VGND sg13g2_fill_1
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_34_159 VPWR VGND sg13g2_decap_8
X_2880_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[0\] _0773_ _0445_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_896 VPWR VGND sg13g2_decap_8
XFILLER_30_310 VPWR VGND sg13g2_fill_2
XFILLER_30_387 VPWR VGND sg13g2_decap_4
X_4550_ _2164_ _2177_ _2141_ _2179_ VPWR VGND sg13g2_nand3_1
X_4481_ _2115_ _2097_ _2114_ VPWR VGND sg13g2_xnor2_1
X_3501_ VGND VPWR _1170_ _1169_ _1148_ sg13g2_or2_1
X_3432_ _1100_ VPWR _1101_ VGND _1094_ _1095_ sg13g2_o21ai_1
X_3363_ _0834_ _0922_ videogen.fancy_shader.video_y\[4\] _1043_ VPWR VGND sg13g2_nand3_1
XFILLER_44_1006 VPWR VGND sg13g2_decap_8
X_5102_ net283 VGND VPWR _0526_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\]
+ _0174_ sg13g2_dfrbpq_1
X_3294_ videogen.fancy_shader.video_y\[1\] videogen.fancy_shader.n646\[1\] _0986_
+ VPWR VGND sg13g2_nor2_1
X_5033_ net178 VGND VPWR _0461_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\]
+ _0118_ sg13g2_dfrbpq_1
XFILLER_25_126 VPWR VGND sg13g2_decap_4
XFILLER_25_137 VPWR VGND sg13g2_decap_8
X_4817_ net691 net741 _0247_ VPWR VGND sg13g2_nor2_1
XFILLER_21_332 VPWR VGND sg13g2_fill_1
XFILLER_22_855 VPWR VGND sg13g2_decap_8
XFILLER_31_26 VPWR VGND sg13g2_fill_1
X_4748_ net673 net725 _0178_ VPWR VGND sg13g2_nor2_1
X_5013__218 VPWR VGND net218 sg13g2_tiehi
X_4679_ net675 net727 _0109_ VPWR VGND sg13g2_nor2_1
Xoutput15 net15 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_16_104 VPWR VGND sg13g2_decap_4
XFILLER_16_148 VPWR VGND sg13g2_fill_1
XFILLER_31_107 VPWR VGND sg13g2_fill_1
XFILLER_12_321 VPWR VGND sg13g2_fill_1
XFILLER_12_332 VPWR VGND sg13g2_fill_1
XFILLER_13_855 VPWR VGND sg13g2_decap_8
XFILLER_8_336 VPWR VGND sg13g2_fill_1
XFILLER_8_369 VPWR VGND sg13g2_decap_8
XFILLER_39_218 VPWR VGND sg13g2_decap_8
XFILLER_36_947 VPWR VGND sg13g2_fill_2
X_4860__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_36_969 VPWR VGND sg13g2_decap_8
XFILLER_35_424 VPWR VGND sg13g2_fill_2
X_3981_ _1645_ _1646_ _1647_ _1648_ _1649_ VPWR VGND sg13g2_nor4_1
X_2932_ _0714_ _0728_ _0785_ VPWR VGND sg13g2_nor2_2
X_2863_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\] net757 _0767_ _0456_
+ VPWR VGND sg13g2_mux2_1
X_2794_ _0728_ _0745_ _0751_ VPWR VGND sg13g2_nor2_2
X_4602_ net662 net714 _0032_ VPWR VGND sg13g2_nor2_1
X_4533_ VGND VPWR _2057_ _2162_ _2163_ net572 sg13g2_a21oi_1
XFILLER_8_870 VPWR VGND sg13g2_decap_8
X_4464_ _2099_ _2096_ _2098_ _2095_ _0863_ VPWR VGND sg13g2_a22oi_1
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
X_3415_ _1084_ videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.n646\[5\]
+ VPWR VGND sg13g2_nand2_1
X_4395_ _2040_ _2037_ _2039_ VPWR VGND sg13g2_xnor2_1
X_3346_ net608 _0922_ _1030_ VPWR VGND sg13g2_and2_1
X_3277_ _0975_ _0808_ _0956_ VPWR VGND sg13g2_nand2_2
X_5016_ net212 VGND VPWR _0444_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\]
+ _0101_ sg13g2_dfrbpq_1
XFILLER_27_903 VPWR VGND sg13g2_fill_1
XFILLER_27_914 VPWR VGND sg13g2_decap_8
X_4881__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_34_490 VPWR VGND sg13g2_fill_2
XFILLER_42_36 VPWR VGND sg13g2_decap_4
XFILLER_21_195 VPWR VGND sg13g2_fill_1
XFILLER_27_1012 VPWR VGND sg13g2_decap_8
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_45_711 VPWR VGND sg13g2_fill_1
XFILLER_45_755 VPWR VGND sg13g2_fill_2
XFILLER_44_221 VPWR VGND sg13g2_fill_1
XFILLER_18_947 VPWR VGND sg13g2_decap_8
XFILLER_33_917 VPWR VGND sg13g2_decap_8
X_5174__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_16_70 VPWR VGND sg13g2_decap_8
XFILLER_9_601 VPWR VGND sg13g2_decap_8
XFILLER_41_972 VPWR VGND sg13g2_decap_8
X_5135__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_34_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_482 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_fill_1
XFILLER_8_166 VPWR VGND sg13g2_decap_8
XFILLER_5_840 VPWR VGND sg13g2_decap_8
XFILLER_5_895 VPWR VGND sg13g2_decap_8
X_4180_ _1842_ _1841_ _1831_ VPWR VGND sg13g2_nand2b_1
X_3200_ _0681_ _0810_ _0923_ _0300_ VPWR VGND sg13g2_nor3_1
X_3131_ _0858_ net599 _0856_ _0861_ VPWR VGND sg13g2_mux2_1
X_3062_ VGND VPWR _0835_ _0845_ net17 _0836_ sg13g2_a21oi_1
XFILLER_24_906 VPWR VGND sg13g2_decap_8
XFILLER_35_298 VPWR VGND sg13g2_fill_1
X_3964_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\] net562 _1632_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_950 VPWR VGND sg13g2_decap_8
X_2915_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\] _0780_ _0417_
+ VPWR VGND sg13g2_mux2_1
X_3895_ net598 _1558_ _1563_ _1564_ VPWR VGND sg13g2_nor3_1
XFILLER_31_471 VPWR VGND sg13g2_decap_8
X_2846_ _0737_ _0758_ _0763_ VPWR VGND sg13g2_nor2_2
XFILLER_31_482 VPWR VGND sg13g2_fill_2
XFILLER_12_39 VPWR VGND sg13g2_fill_2
X_2777_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\] _0747_ _0531_
+ VPWR VGND sg13g2_mux2_1
XFILLER_2_309 VPWR VGND sg13g2_decap_8
X_4516_ _2146_ _2142_ _2144_ VPWR VGND sg13g2_xnor2_1
X_4447_ VGND VPWR _0654_ _2081_ _0619_ _2082_ sg13g2_a21oi_1
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
Xfanout613 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\] net613 VPWR VGND
+ sg13g2_buf_2
Xfanout624 net627 net624 VPWR VGND sg13g2_buf_1
Xfanout635 net640 net635 VPWR VGND sg13g2_buf_8
Xfanout657 net659 net657 VPWR VGND sg13g2_buf_8
X_4378_ _0905_ VPWR _2023_ VGND _0901_ _0902_ sg13g2_o21ai_1
Xfanout646 net648 net646 VPWR VGND sg13g2_buf_8
X_3329_ _0942_ _1018_ _1019_ VPWR VGND sg13g2_nor2b_2
Xfanout679 net681 net679 VPWR VGND sg13g2_buf_8
Xfanout668 net671 net668 VPWR VGND sg13g2_buf_8
XFILLER_46_519 VPWR VGND sg13g2_fill_2
XFILLER_39_560 VPWR VGND sg13g2_decap_4
XFILLER_37_25 VPWR VGND sg13g2_decap_8
XFILLER_27_744 VPWR VGND sg13g2_decap_4
XFILLER_42_703 VPWR VGND sg13g2_decap_4
XFILLER_26_232 VPWR VGND sg13g2_fill_2
XFILLER_42_758 VPWR VGND sg13g2_decap_8
XFILLER_41_257 VPWR VGND sg13g2_fill_2
XFILLER_23_972 VPWR VGND sg13g2_decap_8
XFILLER_2_810 VPWR VGND sg13g2_decap_8
XFILLER_49_302 VPWR VGND sg13g2_decap_8
XFILLER_2_887 VPWR VGND sg13g2_decap_8
XFILLER_40_1020 VPWR VGND sg13g2_decap_8
XFILLER_18_755 VPWR VGND sg13g2_decap_4
XFILLER_18_799 VPWR VGND sg13g2_decap_4
X_4859__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_13_460 VPWR VGND sg13g2_decap_8
XFILLER_14_994 VPWR VGND sg13g2_decap_8
XFILLER_43_90 VPWR VGND sg13g2_decap_4
X_2700_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\] net786 _0725_ _0586_
+ VPWR VGND sg13g2_mux2_1
X_3680_ _1348_ VPWR _1349_ VGND _1312_ _1324_ sg13g2_o21ai_1
X_2631_ _0677_ _0682_ _0684_ VPWR VGND sg13g2_nor2_2
X_4301_ _1962_ _1868_ _1235_ _1963_ VPWR VGND sg13g2_a21o_2
X_4232_ _1894_ _1892_ _1893_ VPWR VGND sg13g2_nand2_1
X_4163_ _1818_ _1815_ _1824_ _1825_ VPWR VGND sg13g2_a21o_1
X_3114_ _0851_ net795 _0822_ VPWR VGND sg13g2_nand2_1
X_4094_ _1705_ _1745_ _1753_ _1759_ VPWR VGND sg13g2_nor3_1
X_3045_ videogen.fancy_shader.video_y\[8\] videogen.fancy_shader.video_y\[7\] _0637_
+ _0832_ VPWR VGND videogen.fancy_shader.video_y\[6\] sg13g2_nand4_1
XFILLER_24_703 VPWR VGND sg13g2_fill_1
X_4996_ net251 VGND VPWR _0424_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\]
+ _0081_ sg13g2_dfrbpq_1
X_3947_ _1614_ VPWR _1615_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\]
+ net577 sg13g2_o21ai_1
XFILLER_20_920 VPWR VGND sg13g2_decap_8
X_3878_ _1543_ _1544_ _1545_ _1546_ _1547_ VPWR VGND sg13g2_nor4_1
X_2829_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[1\] _0759_ _0482_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_997 VPWR VGND sg13g2_decap_8
XFILLER_2_106 VPWR VGND sg13g2_decap_8
XFILLER_2_117 VPWR VGND sg13g2_fill_2
XFILLER_47_806 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_24_1004 VPWR VGND sg13g2_decap_8
XFILLER_27_585 VPWR VGND sg13g2_decap_8
XFILLER_14_235 VPWR VGND sg13g2_fill_1
XFILLER_15_758 VPWR VGND sg13g2_decap_8
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_7_913 VPWR VGND sg13g2_decap_8
XFILLER_6_401 VPWR VGND sg13g2_fill_2
XFILLER_31_1019 VPWR VGND sg13g2_decap_8
XFILLER_6_423 VPWR VGND sg13g2_fill_1
XFILLER_13_82 VPWR VGND sg13g2_fill_1
XFILLER_2_684 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_49_121 VPWR VGND sg13g2_decap_8
XFILLER_49_143 VPWR VGND sg13g2_decap_8
XFILLER_38_839 VPWR VGND sg13g2_decap_8
XFILLER_37_349 VPWR VGND sg13g2_fill_1
X_4850_ net138 VGND VPWR _0278_ red_tmds_par\[7\] net641 sg13g2_dfrbpq_1
X_3801_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[1\] net579 _1470_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_205 VPWR VGND sg13g2_fill_1
XFILLER_14_791 VPWR VGND sg13g2_decap_8
X_4781_ net668 net719 _0211_ VPWR VGND sg13g2_nor2_1
XFILLER_33_599 VPWR VGND sg13g2_fill_1
X_3732_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\] net580 _1401_ VPWR
+ VGND sg13g2_nor2_1
X_3663_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\] net550 _1332_ VPWR
+ VGND sg13g2_nor2_1
X_2614_ VPWR _0669_ net417 VGND sg13g2_inv_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_3594_ VGND VPWR _1263_ _1262_ _1259_ sg13g2_or2_1
X_5195_ net148 VGND VPWR _0619_ tmds_green.dc_balancing_reg\[1\] net645 sg13g2_dfrbpq_2
X_4215_ _1877_ _1089_ _1875_ VPWR VGND sg13g2_xnor2_1
X_4146_ VPWR _1808_ _1807_ VGND sg13g2_inv_1
X_4077_ _1734_ VPWR _1742_ VGND _1738_ _1740_ sg13g2_o21ai_1
X_3028_ VGND VPWR _0824_ videogen.test_lut_thingy.pixel_feeder_inst.state\[3\] videogen.test_lut_thingy.pixel_feeder_inst.state\[1\]
+ sg13g2_or2_1
X_5124__193 VPWR VGND net193 sg13g2_tiehi
X_4979_ net288 VGND VPWR _0407_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\]
+ _0064_ sg13g2_dfrbpq_1
Xclkload3 VPWR clkload3/Y clknet_3_5__leaf_clk_regs VGND sg13g2_inv_1
XFILLER_20_794 VPWR VGND sg13g2_decap_8
XFILLER_19_349 VPWR VGND sg13g2_fill_2
XFILLER_15_511 VPWR VGND sg13g2_fill_2
XFILLER_15_522 VPWR VGND sg13g2_fill_2
XFILLER_42_363 VPWR VGND sg13g2_fill_1
XFILLER_30_503 VPWR VGND sg13g2_decap_4
XFILLER_15_599 VPWR VGND sg13g2_fill_1
XFILLER_7_721 VPWR VGND sg13g2_fill_2
XFILLER_40_80 VPWR VGND sg13g2_decap_8
XFILLER_7_787 VPWR VGND sg13g2_decap_4
X_5110__248 VPWR VGND net248 sg13g2_tiehi
X_4000_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\] net589 _1668_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_27_4 VPWR VGND sg13g2_fill_1
XFILLER_38_647 VPWR VGND sg13g2_decap_8
XFILLER_38_658 VPWR VGND sg13g2_fill_2
X_4902_ net46 VGND VPWR _0330_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\]
+ net630 sg13g2_dfrbpq_1
X_4833_ net650 net702 _0261_ VPWR VGND sg13g2_nor2_1
XFILLER_33_396 VPWR VGND sg13g2_decap_8
X_4764_ net662 net714 _0194_ VPWR VGND sg13g2_nor2_1
X_3715_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\] net589 _1384_ VPWR
+ VGND sg13g2_nor2_1
X_4695_ net680 net730 _0125_ VPWR VGND sg13g2_nor2_1
X_3646_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\] net569 _1315_ VPWR
+ VGND sg13g2_nor2_1
X_3577_ _1138_ _1173_ _1246_ VPWR VGND sg13g2_nor2_1
X_5247_ net801 VGND VPWR serialize.n427\[8\] serialize.n411\[6\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
Xhold15 serialize.n431\[6\] VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold37 serialize.n411\[4\] VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold26 serialize.n411\[7\] VPWR VGND net431 sg13g2_dlygate4sd3_1
XFILLER_29_37 VPWR VGND sg13g2_fill_2
X_5178_ net397 VGND VPWR _0602_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\]
+ _0250_ sg13g2_dfrbpq_1
X_4129_ _1793_ _1495_ _1694_ VPWR VGND sg13g2_nand2_1
XFILLER_45_25 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_fill_2
XFILLER_28_179 VPWR VGND sg13g2_fill_2
XFILLER_25_842 VPWR VGND sg13g2_fill_1
XFILLER_24_352 VPWR VGND sg13g2_decap_8
XFILLER_25_886 VPWR VGND sg13g2_decap_8
XFILLER_24_374 VPWR VGND sg13g2_fill_1
XFILLER_4_702 VPWR VGND sg13g2_fill_1
XFILLER_4_768 VPWR VGND sg13g2_decap_4
XFILLER_10_83 VPWR VGND sg13g2_decap_4
X_5143__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_0_985 VPWR VGND sg13g2_decap_8
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_19_179 VPWR VGND sg13g2_decap_4
XFILLER_35_617 VPWR VGND sg13g2_decap_4
XFILLER_37_1014 VPWR VGND sg13g2_decap_8
X_5138__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_42_182 VPWR VGND sg13g2_decap_8
X_4977__292 VPWR VGND net292 sg13g2_tiehi
X_3500_ _1134_ _1136_ _1146_ _1168_ _1169_ VPWR VGND sg13g2_nor4_1
XFILLER_7_551 VPWR VGND sg13g2_decap_8
X_4480_ _2114_ _2101_ _2112_ VPWR VGND sg13g2_xnor2_1
X_3431_ _1096_ _1099_ _1100_ VPWR VGND sg13g2_and2_1
X_3362_ videogen.fancy_shader.video_y\[4\] _1041_ _1042_ VPWR VGND sg13g2_nor2_1
X_5101_ net287 VGND VPWR _0525_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\]
+ _0173_ sg13g2_dfrbpq_1
XFILLER_39_912 VPWR VGND sg13g2_fill_2
XFILLER_39_901 VPWR VGND sg13g2_fill_2
X_3293_ _0985_ videogen.fancy_shader.video_y\[1\] videogen.fancy_shader.n646\[1\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_400 VPWR VGND sg13g2_fill_1
X_5032_ net180 VGND VPWR _0460_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\]
+ _0117_ sg13g2_dfrbpq_1
XFILLER_38_433 VPWR VGND sg13g2_fill_2
XFILLER_26_617 VPWR VGND sg13g2_decap_8
X_4816_ net688 net740 _0246_ VPWR VGND sg13g2_nor2_1
XFILLER_21_344 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_33_193 VPWR VGND sg13g2_fill_2
XFILLER_21_388 VPWR VGND sg13g2_decap_4
X_4747_ net674 net726 _0177_ VPWR VGND sg13g2_nor2_1
XFILLER_31_38 VPWR VGND sg13g2_decap_8
X_4678_ net675 net727 _0108_ VPWR VGND sg13g2_nor2_1
X_3629_ VGND VPWR _1243_ _1296_ _1298_ _0662_ sg13g2_a21oi_1
Xoutput16 net16 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_738 VPWR VGND sg13g2_decap_8
X_5140__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_16_116 VPWR VGND sg13g2_fill_1
XFILLER_24_171 VPWR VGND sg13g2_decap_4
X_5061__63 VPWR VGND net63 sg13g2_tiehi
XFILLER_4_510 VPWR VGND sg13g2_decap_4
XFILLER_4_543 VPWR VGND sg13g2_fill_2
X_5181__308 VPWR VGND net308 sg13g2_tiehi
XFILLER_0_782 VPWR VGND sg13g2_decap_8
XFILLER_48_775 VPWR VGND sg13g2_decap_4
XFILLER_47_274 VPWR VGND sg13g2_decap_4
XFILLER_36_937 VPWR VGND sg13g2_fill_2
X_3980_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\] net564 _1648_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_44_992 VPWR VGND sg13g2_decap_8
X_2931_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\] _0784_ _0405_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_672 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_15_193 VPWR VGND sg13g2_fill_2
XFILLER_31_653 VPWR VGND sg13g2_fill_1
X_2862_ _0707_ _0758_ _0767_ VPWR VGND sg13g2_nor2_2
X_4601_ net660 net712 _0031_ VPWR VGND sg13g2_nor2_1
XFILLER_30_141 VPWR VGND sg13g2_decap_8
X_2793_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\] net789 _0750_ _0518_
+ VPWR VGND sg13g2_mux2_1
X_4532_ _2162_ _2155_ _2161_ VPWR VGND sg13g2_nand2_1
XFILLER_7_62 VPWR VGND sg13g2_fill_2
XFILLER_7_51 VPWR VGND sg13g2_fill_1
X_4463_ _0863_ _2097_ _2098_ VPWR VGND sg13g2_nor2_1
X_3414_ videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.n646\[5\] _1083_
+ VPWR VGND sg13g2_nor2_1
Xfanout806 rst_n net806 VPWR VGND sg13g2_buf_8
X_4394_ _2039_ tmds_red.dc_balancing_reg\[4\] _2038_ VPWR VGND sg13g2_xnor2_1
X_4869__101 VPWR VGND net101 sg13g2_tiehi
X_3345_ VGND VPWR _0641_ _1028_ _0355_ _1029_ sg13g2_a21oi_1
X_3276_ _0967_ _0974_ _0333_ VPWR VGND sg13g2_nor2_1
X_5015_ net214 VGND VPWR _0443_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\]
+ _0100_ sg13g2_dfrbpq_1
XFILLER_38_285 VPWR VGND sg13g2_fill_2
XFILLER_26_425 VPWR VGND sg13g2_decap_4
XFILLER_21_163 VPWR VGND sg13g2_decap_8
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_1_557 VPWR VGND sg13g2_decap_8
XFILLER_18_926 VPWR VGND sg13g2_decap_8
XFILLER_44_233 VPWR VGND sg13g2_fill_1
XFILLER_17_458 VPWR VGND sg13g2_decap_4
XFILLER_34_1006 VPWR VGND sg13g2_decap_8
XFILLER_40_472 VPWR VGND sg13g2_fill_2
XFILLER_8_156 VPWR VGND sg13g2_fill_1
XFILLER_32_81 VPWR VGND sg13g2_fill_1
XFILLER_5_874 VPWR VGND sg13g2_decap_8
X_3130_ _0860_ net601 _0856_ VPWR VGND sg13g2_nand2_1
XFILLER_36_712 VPWR VGND sg13g2_decap_4
X_3061_ _0845_ _0843_ _0844_ VPWR VGND sg13g2_nand2_1
XFILLER_35_200 VPWR VGND sg13g2_decap_4
XFILLER_16_480 VPWR VGND sg13g2_fill_2
X_3963_ net620 VPWR _1631_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\]
+ net574 sg13g2_o21ai_1
X_2914_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\] _0780_ _0418_
+ VPWR VGND sg13g2_mux2_1
X_3894_ net618 _1559_ _1560_ _1562_ _1563_ VPWR VGND sg13g2_nor4_1
XFILLER_31_450 VPWR VGND sg13g2_fill_1
X_2845_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\] _0762_ _0469_
+ VPWR VGND sg13g2_mux2_1
X_2776_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\] _0747_ _0532_
+ VPWR VGND sg13g2_mux2_1
X_4515_ _2142_ _2144_ _2145_ VPWR VGND sg13g2_nor2_1
X_4446_ _0852_ VPWR _2082_ VGND _0654_ _2081_ sg13g2_o21ai_1
Xfanout603 net604 net603 VPWR VGND sg13g2_buf_2
Xfanout614 net615 net614 VPWR VGND sg13g2_buf_8
X_4377_ _2005_ VPWR _2022_ VGND _1999_ _2003_ sg13g2_o21ai_1
X_3328_ _1009_ _1017_ _1018_ VPWR VGND sg13g2_nor2b_2
Xfanout658 net659 net658 VPWR VGND sg13g2_buf_1
Xfanout636 net640 net636 VPWR VGND sg13g2_buf_8
Xfanout647 net648 net647 VPWR VGND sg13g2_buf_8
Xfanout625 net627 net625 VPWR VGND sg13g2_buf_8
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
XFILLER_37_48 VPWR VGND sg13g2_decap_8
X_3259_ _0809_ _0962_ _0963_ _0327_ VPWR VGND sg13g2_nor3_1
XFILLER_39_594 VPWR VGND sg13g2_fill_1
XFILLER_42_737 VPWR VGND sg13g2_fill_1
XFILLER_14_439 VPWR VGND sg13g2_fill_2
XFILLER_23_951 VPWR VGND sg13g2_decap_8
XFILLER_22_450 VPWR VGND sg13g2_fill_1
XFILLER_5_115 VPWR VGND sg13g2_decap_8
XFILLER_5_104 VPWR VGND sg13g2_fill_2
XFILLER_2_866 VPWR VGND sg13g2_decap_8
XFILLER_18_712 VPWR VGND sg13g2_decap_8
XFILLER_17_233 VPWR VGND sg13g2_fill_2
XFILLER_33_704 VPWR VGND sg13g2_decap_8
XFILLER_33_715 VPWR VGND sg13g2_fill_2
XFILLER_17_299 VPWR VGND sg13g2_fill_1
XFILLER_32_247 VPWR VGND sg13g2_decap_4
XFILLER_14_973 VPWR VGND sg13g2_decap_8
XFILLER_32_258 VPWR VGND sg13g2_fill_1
XFILLER_13_494 VPWR VGND sg13g2_fill_1
X_2630_ _0683_ _0682_ VPWR VGND sg13g2_inv_2
X_4300_ _1960_ VPWR _1962_ VGND _1957_ _1958_ sg13g2_o21ai_1
XFILLER_4_192 VPWR VGND sg13g2_decap_4
XFILLER_4_52 VPWR VGND sg13g2_decap_8
X_4231_ VGND VPWR _1893_ _1886_ _1884_ sg13g2_or2_1
X_4913__396 VPWR VGND net396 sg13g2_tiehi
XFILLER_4_63 VPWR VGND sg13g2_fill_2
X_4162_ VGND VPWR _1810_ _1813_ _1824_ _1807_ sg13g2_a21oi_1
X_5083__367 VPWR VGND net367 sg13g2_tiehi
X_3113_ VPWR clk_video _0006_ VGND sg13g2_inv_1
X_4093_ _1745_ _1754_ _1757_ _1758_ VPWR VGND sg13g2_nor3_1
X_3044_ _0831_ videogen.fancy_shader.video_y\[1\] net608 VPWR VGND sg13g2_nand2_1
XFILLER_24_737 VPWR VGND sg13g2_decap_8
XFILLER_36_586 VPWR VGND sg13g2_decap_8
XFILLER_36_597 VPWR VGND sg13g2_fill_1
X_4995_ net253 VGND VPWR _0423_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\]
+ _0080_ sg13g2_dfrbpq_1
XFILLER_23_225 VPWR VGND sg13g2_decap_4
XFILLER_11_409 VPWR VGND sg13g2_fill_2
X_3946_ _1614_ net593 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
X_3877_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\] net562 _1546_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_976 VPWR VGND sg13g2_decap_8
X_2828_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[2\] _0759_ _0483_
+ VPWR VGND sg13g2_mux2_1
X_2759_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\] net777 _0741_ _0543_
+ VPWR VGND sg13g2_mux2_1
X_4429_ _2068_ _2069_ _0612_ VPWR VGND sg13g2_nor2_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_39_391 VPWR VGND sg13g2_fill_1
XFILLER_14_214 VPWR VGND sg13g2_decap_8
XFILLER_15_748 VPWR VGND sg13g2_decap_4
XFILLER_11_910 VPWR VGND sg13g2_decap_8
X_5171__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_10_453 VPWR VGND sg13g2_decap_8
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_13_61 VPWR VGND sg13g2_decap_8
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_1_195 VPWR VGND sg13g2_fill_1
XFILLER_37_306 VPWR VGND sg13g2_fill_2
XFILLER_49_199 VPWR VGND sg13g2_decap_8
XFILLER_18_553 VPWR VGND sg13g2_fill_2
XFILLER_46_895 VPWR VGND sg13g2_decap_8
X_3800_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\] net557 _1469_ VPWR
+ VGND sg13g2_nor2_1
X_4780_ net668 net719 _0210_ VPWR VGND sg13g2_nor2_1
X_3731_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\] net591 _1400_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_228 VPWR VGND sg13g2_decap_8
X_3662_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\] net585 _1331_ VPWR
+ VGND sg13g2_nor2_1
X_2613_ VPWR _0668_ net414 VGND sg13g2_inv_1
X_3593_ net544 _1257_ _1262_ VPWR VGND sg13g2_nor2_1
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_5_490 VPWR VGND sg13g2_decap_8
X_4987__272 VPWR VGND net272 sg13g2_tiehi
X_5194_ net163 VGND VPWR _0618_ blue_tmds_par\[9\] net637 sg13g2_dfrbpq_1
X_4214_ _1073_ _1086_ _1087_ _1876_ VGND VPWR _1870_ sg13g2_nor4_2
X_4145_ _1807_ _1713_ _1806_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_862 VPWR VGND sg13g2_fill_2
X_4076_ _1738_ _1740_ _1741_ VPWR VGND sg13g2_nor2_1
X_3027_ _0823_ videogen.test_lut_thingy.pixel_feeder_inst.state\[1\] _0807_ VPWR VGND
+ sg13g2_nand2b_1
XFILLER_24_501 VPWR VGND sg13g2_fill_2
X_4978_ net290 VGND VPWR _0406_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\]
+ _0063_ sg13g2_dfrbpq_1
X_3929_ net626 VPWR _1597_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\]
+ net581 sg13g2_o21ai_1
Xclkload4 VPWR clkload4/Y clknet_3_7__leaf_clk_regs VGND sg13g2_inv_1
XFILLER_4_939 VPWR VGND sg13g2_decap_8
XFILLER_3_405 VPWR VGND sg13g2_fill_2
X_5131__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
XFILLER_42_331 VPWR VGND sg13g2_decap_4
XFILLER_42_375 VPWR VGND sg13g2_fill_2
XFILLER_24_71 VPWR VGND sg13g2_decap_8
XFILLER_24_93 VPWR VGND sg13g2_decap_8
XFILLER_30_548 VPWR VGND sg13g2_fill_2
XFILLER_30_559 VPWR VGND sg13g2_decap_8
XFILLER_11_773 VPWR VGND sg13g2_fill_2
XFILLER_7_755 VPWR VGND sg13g2_fill_1
XFILLER_6_232 VPWR VGND sg13g2_fill_2
XFILLER_7_799 VPWR VGND sg13g2_decap_8
XFILLER_40_92 VPWR VGND sg13g2_fill_2
XFILLER_41_7 VPWR VGND sg13g2_fill_2
XFILLER_3_983 VPWR VGND sg13g2_decap_8
XFILLER_19_862 VPWR VGND sg13g2_decap_8
XFILLER_45_180 VPWR VGND sg13g2_decap_4
X_4901_ net48 VGND VPWR _0329_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\]
+ net648 sg13g2_dfrbpq_2
XFILLER_21_504 VPWR VGND sg13g2_decap_8
X_4832_ net650 net702 _0260_ VPWR VGND sg13g2_nor2_1
XFILLER_14_1015 VPWR VGND sg13g2_decap_8
X_4763_ net668 net719 _0193_ VPWR VGND sg13g2_nor2_1
X_3714_ net616 VPWR _1383_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[2\]
+ net579 sg13g2_o21ai_1
X_4694_ net679 net731 _0124_ VPWR VGND sg13g2_nor2_1
X_3645_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\] net558 _1314_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_18 VPWR VGND sg13g2_fill_2
X_3576_ _1220_ VPWR _1245_ VGND _1063_ _1231_ sg13g2_o21ai_1
XFILLER_0_408 VPWR VGND sg13g2_fill_2
X_5246_ net802 VGND VPWR serialize.n427\[7\] serialize.n411\[5\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
Xhold38 serialize.n417\[4\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold16 serialize.n411\[0\] VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold27 clockdiv.q0 VPWR VGND net432 sg13g2_dlygate4sd3_1
X_5177_ net41 VGND VPWR _0601_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\]
+ _0249_ sg13g2_dfrbpq_1
XFILLER_28_136 VPWR VGND sg13g2_decap_8
XFILLER_29_648 VPWR VGND sg13g2_decap_4
X_4128_ _0377_ _1790_ _1792_ VPWR VGND sg13g2_nand2_1
XFILLER_29_659 VPWR VGND sg13g2_fill_1
X_4059_ _1718_ _1719_ _1721_ _1722_ _1724_ VPWR VGND sg13g2_nor4_1
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_24_342 VPWR VGND sg13g2_fill_1
XFILLER_25_865 VPWR VGND sg13g2_decap_8
XFILLER_40_835 VPWR VGND sg13g2_fill_1
Xclkbuf_regs_0_clk clk clk_regs VPWR VGND sg13g2_buf_8
XFILLER_0_964 VPWR VGND sg13g2_decap_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_fill_2
XFILLER_19_125 VPWR VGND sg13g2_decap_4
XFILLER_15_320 VPWR VGND sg13g2_fill_2
XFILLER_16_821 VPWR VGND sg13g2_fill_1
XFILLER_27_180 VPWR VGND sg13g2_decap_8
XFILLER_30_312 VPWR VGND sg13g2_fill_1
X_3430_ videogen.fancy_shader.n646\[6\] videogen.fancy_shader.video_y\[6\] _1099_
+ VPWR VGND sg13g2_xor2_1
X_3361_ net750 _1040_ _1041_ _0359_ VPWR VGND sg13g2_nor3_1
X_5100_ net291 VGND VPWR _0524_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\]
+ _0172_ sg13g2_dfrbpq_1
X_5031_ net182 VGND VPWR _0459_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\]
+ _0116_ sg13g2_dfrbpq_1
X_3292_ VGND VPWR videogen.fancy_shader.n646\[1\] _0981_ _0984_ videogen.fancy_shader.n646\[2\]
+ sg13g2_a21oi_1
XFILLER_39_946 VPWR VGND sg13g2_fill_2
X_4893__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_38_445 VPWR VGND sg13g2_fill_1
XFILLER_25_106 VPWR VGND sg13g2_fill_2
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_34_640 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_fill_1
XFILLER_22_824 VPWR VGND sg13g2_decap_8
X_4815_ net688 net740 _0245_ VPWR VGND sg13g2_nor2_1
XFILLER_31_17 VPWR VGND sg13g2_decap_8
X_4839__153 VPWR VGND net153 sg13g2_tiehi
X_4746_ net673 net725 _0176_ VPWR VGND sg13g2_nor2_1
X_4677_ net687 net735 _0107_ VPWR VGND sg13g2_nor2_1
X_3628_ net750 _0662_ _1297_ VPWR VGND sg13g2_nor2_1
Xoutput17 net17 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_227 VPWR VGND sg13g2_fill_2
XFILLER_0_205 VPWR VGND sg13g2_decap_4
X_3559_ VGND VPWR _1215_ _1217_ _1228_ _1211_ sg13g2_a21oi_1
X_5229_ net799 VGND VPWR net434 serialize.n417\[1\] clknet_3_2__leaf_clk_regs sg13g2_dfrbpq_1
XFILLER_48_209 VPWR VGND sg13g2_fill_2
XFILLER_45_949 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_fill_1
XFILLER_44_437 VPWR VGND sg13g2_fill_2
XFILLER_16_139 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_25_684 VPWR VGND sg13g2_decap_8
XFILLER_12_345 VPWR VGND sg13g2_fill_2
XFILLER_9_839 VPWR VGND sg13g2_decap_8
XFILLER_12_367 VPWR VGND sg13g2_decap_8
XFILLER_8_349 VPWR VGND sg13g2_decap_4
XFILLER_21_83 VPWR VGND sg13g2_fill_2
XFILLER_0_761 VPWR VGND sg13g2_decap_8
XFILLER_36_905 VPWR VGND sg13g2_fill_2
XFILLER_35_437 VPWR VGND sg13g2_decap_8
XFILLER_35_448 VPWR VGND sg13g2_fill_1
XFILLER_44_971 VPWR VGND sg13g2_decap_8
X_2930_ net776 videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\] _0784_ _0406_
+ VPWR VGND sg13g2_mux2_1
XFILLER_22_109 VPWR VGND sg13g2_fill_1
XFILLER_43_492 VPWR VGND sg13g2_decap_4
X_4600_ net660 net712 _0030_ VPWR VGND sg13g2_nor2_1
X_2861_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\] _0766_ _0457_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_665 VPWR VGND sg13g2_decap_8
XFILLER_8_850 VPWR VGND sg13g2_fill_2
X_2792_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\] net779 _0750_ _0519_
+ VPWR VGND sg13g2_mux2_1
X_5190__195 VPWR VGND net195 sg13g2_tiehi
X_4531_ _2161_ _2149_ net602 VPWR VGND sg13g2_nand2b_1
X_4462_ VGND VPWR _2090_ _2097_ _0652_ net599 sg13g2_a21oi_2
XFILLER_7_96 VPWR VGND sg13g2_decap_8
X_5012__220 VPWR VGND net220 sg13g2_tiehi
X_3413_ _1082_ _1080_ _1081_ VPWR VGND sg13g2_xnor2_1
X_4393_ VGND VPWR _0666_ _2023_ _2038_ _0902_ sg13g2_a21oi_1
X_3344_ net795 VPWR _1029_ VGND _0641_ _1028_ sg13g2_o21ai_1
X_3275_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] _0973_ _0974_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_39_721 VPWR VGND sg13g2_fill_1
X_5014_ net216 VGND VPWR _0442_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\]
+ _0099_ sg13g2_dfrbpq_1
X_5162__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_38_264 VPWR VGND sg13g2_decap_8
XFILLER_27_949 VPWR VGND sg13g2_decap_8
X_4923__376 VPWR VGND net376 sg13g2_tiehi
XFILLER_22_621 VPWR VGND sg13g2_fill_1
XFILLER_34_492 VPWR VGND sg13g2_fill_1
XFILLER_10_816 VPWR VGND sg13g2_fill_2
X_4729_ net649 net701 _0159_ VPWR VGND sg13g2_nor2_1
XFILLER_1_536 VPWR VGND sg13g2_decap_8
XFILLER_18_905 VPWR VGND sg13g2_decap_8
XFILLER_29_242 VPWR VGND sg13g2_fill_1
XFILLER_45_746 VPWR VGND sg13g2_fill_1
XFILLER_44_245 VPWR VGND sg13g2_fill_1
XFILLER_26_993 VPWR VGND sg13g2_decap_8
XFILLER_40_451 VPWR VGND sg13g2_decap_8
XFILLER_8_135 VPWR VGND sg13g2_fill_1
XFILLER_9_658 VPWR VGND sg13g2_fill_1
XFILLER_13_698 VPWR VGND sg13g2_fill_2
X_5185__242 VPWR VGND net242 sg13g2_tiehi
X_3060_ _0840_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\]
+ _0844_ VPWR VGND sg13g2_a21o_1
XFILLER_48_573 VPWR VGND sg13g2_decap_4
XFILLER_35_223 VPWR VGND sg13g2_fill_1
XFILLER_17_982 VPWR VGND sg13g2_decap_8
X_3962_ net598 _1624_ _1629_ _1630_ VPWR VGND sg13g2_nor3_1
X_2913_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\] _0780_ _0419_
+ VPWR VGND sg13g2_mux2_1
X_3893_ _1561_ VPWR _1562_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\]
+ net561 sg13g2_o21ai_1
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_2844_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\] _0762_ _0470_
+ VPWR VGND sg13g2_mux2_1
X_2775_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\] _0747_ _0533_
+ VPWR VGND sg13g2_mux2_1
X_4514_ _2143_ VPWR _2144_ VGND tmds_blue.dc_balancing_reg\[1\] _2139_ sg13g2_o21ai_1
X_4836__156 VPWR VGND net156 sg13g2_tiehi
X_4445_ _2079_ _2080_ _2081_ VPWR VGND sg13g2_nor2_2
Xfanout615 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net615 VPWR VGND
+ sg13g2_buf_8
Xfanout604 tmds_blue.n100 net604 VPWR VGND sg13g2_buf_1
X_4376_ VGND VPWR _2016_ _2021_ _0511_ net571 sg13g2_a21oi_1
Xfanout637 net638 net637 VPWR VGND sg13g2_buf_8
Xfanout648 clk_video net648 VPWR VGND sg13g2_buf_8
X_3327_ _1016_ _1013_ _1017_ VPWR VGND sg13g2_nor2b_1
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_1
Xfanout659 net672 net659 VPWR VGND sg13g2_buf_2
X_3258_ net596 _0646_ net578 _0956_ _0963_ VPWR VGND sg13g2_nor4_1
X_5127__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
X_3189_ _0916_ VPWR _0917_ VGND net547 _0912_ sg13g2_o21ai_1
XFILLER_15_919 VPWR VGND sg13g2_decap_8
XFILLER_14_429 VPWR VGND sg13g2_fill_1
XFILLER_23_930 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_fill_1
XFILLER_10_635 VPWR VGND sg13g2_decap_8
XFILLER_10_646 VPWR VGND sg13g2_fill_1
XFILLER_10_679 VPWR VGND sg13g2_fill_1
XFILLER_2_845 VPWR VGND sg13g2_decap_8
XFILLER_14_952 VPWR VGND sg13g2_decap_8
X_5113__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_5_672 VPWR VGND sg13g2_fill_2
X_4230_ _1886_ _1891_ _1884_ _1892_ VPWR VGND sg13g2_nand3_1
XFILLER_4_86 VPWR VGND sg13g2_decap_4
X_4161_ _1816_ _1820_ _1821_ _1823_ VPWR VGND sg13g2_or3_1
X_3112_ net677 net729 _0006_ VPWR VGND sg13g2_nor2_1
X_4092_ _1755_ _1756_ _1757_ VPWR VGND sg13g2_and2_1
XFILLER_49_882 VPWR VGND sg13g2_decap_8
X_3043_ _0830_ videogen.fancy_shader.video_y\[4\] videogen.fancy_shader.video_y\[5\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_36_521 VPWR VGND sg13g2_decap_8
X_4994_ net255 VGND VPWR _0422_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\]
+ _0079_ sg13g2_dfrbpq_1
XFILLER_17_1024 VPWR VGND sg13g2_decap_4
X_3945_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\] net564 _1613_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_771 VPWR VGND sg13g2_fill_2
X_3876_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\] net551 _1545_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_955 VPWR VGND sg13g2_decap_8
XFILLER_31_281 VPWR VGND sg13g2_decap_8
X_4906__38 VPWR VGND net38 sg13g2_tiehi
X_2827_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\] _0759_ _0484_
+ VPWR VGND sg13g2_mux2_1
X_2758_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\] net771 _0741_ _0544_
+ VPWR VGND sg13g2_mux2_1
X_4428_ net799 VPWR _2069_ VGND net605 _0667_ sg13g2_o21ai_1
X_2689_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\] _0723_ _0595_
+ VPWR VGND sg13g2_mux2_1
X_4359_ VGND VPWR _2005_ _2004_ _1996_ sg13g2_or2_1
XFILLER_39_370 VPWR VGND sg13g2_decap_8
XFILLER_23_771 VPWR VGND sg13g2_decap_8
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_13_51 VPWR VGND sg13g2_decap_4
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_6_414 VPWR VGND sg13g2_decap_4
XFILLER_10_476 VPWR VGND sg13g2_fill_2
XFILLER_49_178 VPWR VGND sg13g2_decap_8
XFILLER_38_81 VPWR VGND sg13g2_decap_8
XFILLER_18_521 VPWR VGND sg13g2_decap_8
XFILLER_46_874 VPWR VGND sg13g2_decap_8
XFILLER_45_362 VPWR VGND sg13g2_fill_2
XFILLER_33_524 VPWR VGND sg13g2_decap_8
XFILLER_33_557 VPWR VGND sg13g2_decap_8
X_3730_ VPWR _1399_ _1398_ VGND sg13g2_inv_1
X_3661_ net614 VPWR _1330_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\]
+ net561 sg13g2_o21ai_1
X_3592_ VGND VPWR _1255_ _1260_ _1261_ _1253_ sg13g2_a21oi_1
XFILLER_6_970 VPWR VGND sg13g2_decap_8
X_5193_ net171 VGND VPWR _0617_ blue_tmds_par\[8\] net637 sg13g2_dfrbpq_1
X_4213_ _1875_ _1018_ _1874_ VPWR VGND sg13g2_xnor2_1
X_4144_ _1082_ _1121_ _1018_ _1806_ VPWR VGND sg13g2_nand3_1
X_4075_ _1740_ _1707_ _1728_ _1739_ VPWR VGND sg13g2_and3_1
X_3026_ _0822_ _0818_ _0821_ _0817_ _0816_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_513 VPWR VGND sg13g2_fill_2
XFILLER_12_719 VPWR VGND sg13g2_fill_1
X_4977_ net292 VGND VPWR _0405_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\]
+ _0062_ sg13g2_dfrbpq_1
XFILLER_11_207 VPWR VGND sg13g2_fill_2
X_4994__255 VPWR VGND net255 sg13g2_tiehi
XFILLER_20_752 VPWR VGND sg13g2_fill_1
X_3928_ VPWR _0372_ _1596_ VGND sg13g2_inv_1
X_3859_ net624 VPWR _1528_ VGND _1525_ _1527_ sg13g2_o21ai_1
XFILLER_4_918 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
X_4966__313 VPWR VGND net313 sg13g2_tiehi
XFILLER_47_627 VPWR VGND sg13g2_fill_2
X_5103__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_15_513 VPWR VGND sg13g2_fill_1
XFILLER_42_354 VPWR VGND sg13g2_decap_8
XFILLER_11_763 VPWR VGND sg13g2_decap_8
XFILLER_11_796 VPWR VGND sg13g2_decap_4
XFILLER_6_266 VPWR VGND sg13g2_fill_2
XFILLER_3_962 VPWR VGND sg13g2_decap_8
XFILLER_2_472 VPWR VGND sg13g2_decap_4
XFILLER_34_7 VPWR VGND sg13g2_fill_2
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_38_616 VPWR VGND sg13g2_fill_2
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_fill_1
XFILLER_1_65 VPWR VGND sg13g2_fill_1
XFILLER_19_830 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_fill_2
X_4900_ net50 VGND VPWR _0328_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[4\]
+ net630 sg13g2_dfrbpq_2
X_4831_ net650 net702 _0259_ VPWR VGND sg13g2_nor2_1
XFILLER_33_365 VPWR VGND sg13g2_decap_4
X_5193__171 VPWR VGND net171 sg13g2_tiehi
X_4762_ net669 net719 _0192_ VPWR VGND sg13g2_nor2_1
XFILLER_21_549 VPWR VGND sg13g2_decap_8
X_3713_ _0646_ _1376_ _1381_ _1382_ VPWR VGND sg13g2_nor3_1
X_4693_ net679 net731 _0123_ VPWR VGND sg13g2_nor2_1
X_3644_ net597 VPWR _1313_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\]
+ net591 sg13g2_o21ai_1
X_3575_ VPWR VGND _1241_ _1232_ _1240_ _1233_ _1244_ _1234_ sg13g2_a221oi_1
X_5245_ net802 VGND VPWR serialize.n427\[6\] serialize.n411\[4\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
Xhold28 serialize.n417\[3\] VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold17 serialize.n411\[2\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold39 serialize.n429\[4\] VPWR VGND net444 sg13g2_dlygate4sd3_1
X_5176_ net57 VGND VPWR _0600_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\]
+ _0248_ sg13g2_dfrbpq_1
XFILLER_29_605 VPWR VGND sg13g2_fill_2
X_4127_ _1591_ _1398_ _1791_ _1792_ VPWR VGND sg13g2_a21o_1
X_4058_ _1721_ _1722_ _1723_ VPWR VGND sg13g2_nor2_2
X_5022__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_45_49 VPWR VGND sg13g2_decap_8
X_3009_ videogen.fancy_shader.video_x\[8\] videogen.fancy_shader.video_x\[9\] _0806_
+ VPWR VGND sg13g2_and2_1
XFILLER_24_321 VPWR VGND sg13g2_decap_8
XFILLER_24_398 VPWR VGND sg13g2_decap_8
XFILLER_4_737 VPWR VGND sg13g2_decap_8
X_4933__356 VPWR VGND net356 sg13g2_tiehi
XFILLER_0_943 VPWR VGND sg13g2_decap_8
XFILLER_48_914 VPWR VGND sg13g2_decap_8
XFILLER_47_446 VPWR VGND sg13g2_decap_8
XFILLER_19_72 VPWR VGND sg13g2_decap_8
XFILLER_47_457 VPWR VGND sg13g2_fill_1
XFILLER_16_844 VPWR VGND sg13g2_fill_1
XFILLER_15_343 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_fill_1
XFILLER_31_847 VPWR VGND sg13g2_fill_1
XFILLER_30_357 VPWR VGND sg13g2_decap_4
X_3360_ _0829_ _1033_ _1041_ VPWR VGND sg13g2_nor2_1
XFILLER_39_903 VPWR VGND sg13g2_fill_1
XFILLER_2_291 VPWR VGND sg13g2_fill_1
X_5030_ net184 VGND VPWR _0458_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\]
+ _0115_ sg13g2_dfrbpq_1
X_3291_ VGND VPWR videogen.fancy_shader.n646\[1\] _0981_ _0347_ _0983_ sg13g2_a21oi_1
XFILLER_34_663 VPWR VGND sg13g2_decap_8
X_5070__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_22_869 VPWR VGND sg13g2_fill_2
X_4814_ net688 net740 _0244_ VPWR VGND sg13g2_nor2_1
X_4745_ net659 net708 _0175_ VPWR VGND sg13g2_nor2_1
X_4676_ net687 net735 _0106_ VPWR VGND sg13g2_nor2_1
X_3627_ _1239_ _1244_ _1294_ _1295_ _1296_ VPWR VGND sg13g2_nor4_1
Xoutput18 net18 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_707 VPWR VGND sg13g2_fill_1
X_3558_ _1222_ VPWR _1227_ VGND _1224_ _1225_ sg13g2_o21ai_1
X_3489_ _1156_ _1157_ _1158_ VPWR VGND sg13g2_nor2_2
XFILLER_0_239 VPWR VGND sg13g2_decap_8
X_5228_ net799 VGND VPWR serialize.n429\[2\] serialize.n417\[0\] clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
X_5159_ net254 VGND VPWR _0583_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[1\]
+ _0231_ sg13g2_dfrbpq_1
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_17_619 VPWR VGND sg13g2_decap_8
XFILLER_40_611 VPWR VGND sg13g2_fill_2
XFILLER_25_663 VPWR VGND sg13g2_fill_1
XFILLER_40_633 VPWR VGND sg13g2_fill_2
XFILLER_13_869 VPWR VGND sg13g2_fill_2
XFILLER_8_306 VPWR VGND sg13g2_decap_8
XFILLER_4_545 VPWR VGND sg13g2_fill_1
XFILLER_0_740 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_fill_2
X_5109__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_36_939 VPWR VGND sg13g2_fill_1
XFILLER_46_81 VPWR VGND sg13g2_decap_8
XFILLER_44_950 VPWR VGND sg13g2_decap_8
XFILLER_15_195 VPWR VGND sg13g2_fill_1
X_2860_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[1\] _0766_ _0458_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_677 VPWR VGND sg13g2_decap_8
X_2791_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\] net768 _0750_ _0520_
+ VPWR VGND sg13g2_mux2_1
XFILLER_12_891 VPWR VGND sg13g2_decap_8
XFILLER_30_176 VPWR VGND sg13g2_decap_8
XFILLER_31_699 VPWR VGND sg13g2_decap_8
X_4530_ VPWR VGND _2155_ _2057_ _2159_ _2060_ _2160_ _2158_ sg13g2_a221oi_1
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
X_4461_ _2096_ _2090_ _2078_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_884 VPWR VGND sg13g2_decap_8
XFILLER_7_372 VPWR VGND sg13g2_decap_8
XFILLER_7_75 VPWR VGND sg13g2_decap_8
X_3412_ _0998_ VPWR _1081_ VGND _0999_ _1008_ sg13g2_o21ai_1
X_4392_ VGND VPWR _2024_ _2032_ _2037_ _2034_ sg13g2_a21oi_1
X_3343_ _0354_ net795 _1027_ _1028_ VPWR VGND sg13g2_and3_1
X_3274_ _0967_ _0972_ _0973_ _0332_ VPWR VGND sg13g2_nor3_1
XFILLER_38_221 VPWR VGND sg13g2_fill_1
XFILLER_38_210 VPWR VGND sg13g2_fill_1
X_5013_ net218 VGND VPWR _0441_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[0\]
+ _0098_ sg13g2_dfrbpq_1
XFILLER_39_777 VPWR VGND sg13g2_decap_8
XFILLER_38_243 VPWR VGND sg13g2_decap_8
XFILLER_27_928 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_fill_2
XFILLER_41_408 VPWR VGND sg13g2_decap_8
XFILLER_22_600 VPWR VGND sg13g2_decap_8
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_21_121 VPWR VGND sg13g2_decap_8
XFILLER_21_143 VPWR VGND sg13g2_decap_8
X_2989_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\] _0800_ _0289_
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_187 VPWR VGND sg13g2_decap_4
X_4728_ net649 net701 _0158_ VPWR VGND sg13g2_nor2_1
XFILLER_5_309 VPWR VGND sg13g2_fill_1
X_4659_ net670 net721 _0089_ VPWR VGND sg13g2_nor2_1
XFILLER_1_515 VPWR VGND sg13g2_decap_8
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_44_213 VPWR VGND sg13g2_decap_4
XFILLER_29_276 VPWR VGND sg13g2_decap_4
XFILLER_26_972 VPWR VGND sg13g2_decap_8
XFILLER_32_408 VPWR VGND sg13g2_fill_2
XFILLER_41_986 VPWR VGND sg13g2_decap_8
XFILLER_13_677 VPWR VGND sg13g2_decap_8
XFILLER_40_496 VPWR VGND sg13g2_decap_8
XFILLER_9_637 VPWR VGND sg13g2_decap_8
XFILLER_13_688 VPWR VGND sg13g2_fill_2
XFILLER_32_94 VPWR VGND sg13g2_fill_1
XFILLER_4_331 VPWR VGND sg13g2_fill_1
XFILLER_48_552 VPWR VGND sg13g2_decap_8
X_3961_ _1625_ _1626_ _1627_ _1628_ _1629_ VPWR VGND sg13g2_nor4_1
XFILLER_17_961 VPWR VGND sg13g2_decap_8
XFILLER_23_408 VPWR VGND sg13g2_fill_1
X_2912_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\] _0780_ _0420_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_482 VPWR VGND sg13g2_fill_1
X_3892_ _1561_ net593 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_31_441 VPWR VGND sg13g2_decap_8
XFILLER_32_964 VPWR VGND sg13g2_decap_8
X_2843_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\] _0762_ _0471_
+ VPWR VGND sg13g2_mux2_1
X_2774_ _0747_ _0722_ _0744_ VPWR VGND sg13g2_nand2_2
X_4513_ _2143_ _2139_ _2138_ VPWR VGND sg13g2_nand2b_1
X_4444_ VGND VPWR _2077_ _2078_ _2080_ net600 sg13g2_a21oi_1
Xfanout605 net607 net605 VPWR VGND sg13g2_buf_8
X_4375_ _2010_ _2020_ _2021_ VPWR VGND sg13g2_nor2_1
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_1
Xfanout649 net651 net649 VPWR VGND sg13g2_buf_8
X_3326_ _1016_ _1014_ _1015_ VPWR VGND sg13g2_xnor2_1
Xfanout616 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net616 VPWR VGND
+ sg13g2_buf_8
Xfanout627 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\] net627 VPWR VGND
+ sg13g2_buf_8
XFILLER_37_39 VPWR VGND sg13g2_decap_4
X_3257_ VGND VPWR net623 _0959_ _0962_ net616 sg13g2_a21oi_1
XFILLER_39_585 VPWR VGND sg13g2_decap_8
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
XFILLER_26_202 VPWR VGND sg13g2_fill_2
X_3188_ _0916_ net547 _0910_ VPWR VGND sg13g2_nand2_1
XFILLER_26_257 VPWR VGND sg13g2_fill_1
XFILLER_23_986 VPWR VGND sg13g2_decap_8
XFILLER_6_618 VPWR VGND sg13g2_decap_8
XFILLER_6_629 VPWR VGND sg13g2_fill_1
XFILLER_5_106 VPWR VGND sg13g2_fill_1
XFILLER_5_139 VPWR VGND sg13g2_fill_2
XFILLER_2_824 VPWR VGND sg13g2_decap_8
X_5030__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_49_316 VPWR VGND sg13g2_decap_4
XFILLER_45_544 VPWR VGND sg13g2_decap_8
XFILLER_17_235 VPWR VGND sg13g2_fill_1
XFILLER_17_257 VPWR VGND sg13g2_decap_8
XFILLER_27_94 VPWR VGND sg13g2_fill_1
XFILLER_32_205 VPWR VGND sg13g2_decap_8
XFILLER_14_931 VPWR VGND sg13g2_decap_8
XFILLER_25_290 VPWR VGND sg13g2_decap_8
XFILLER_13_474 VPWR VGND sg13g2_fill_1
XFILLER_13_485 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_fill_2
XFILLER_4_183 VPWR VGND sg13g2_decap_4
X_4160_ _1816_ _1818_ _1819_ _1821_ _1822_ VPWR VGND sg13g2_nor4_1
XFILLER_4_76 VPWR VGND sg13g2_decap_4
X_3111_ red_tmds_par\[9\] net695 serialize.n427\[9\] VPWR VGND sg13g2_and2_1
XFILLER_49_861 VPWR VGND sg13g2_decap_8
X_4091_ _1756_ _0990_ _1066_ VPWR VGND sg13g2_nand2_1
XFILLER_48_360 VPWR VGND sg13g2_fill_2
X_3042_ _0829_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_36_544 VPWR VGND sg13g2_fill_2
XFILLER_36_555 VPWR VGND sg13g2_decap_8
X_4993_ net257 VGND VPWR _0421_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\]
+ _0078_ sg13g2_dfrbpq_1
XFILLER_17_1003 VPWR VGND sg13g2_decap_8
X_3944_ _1608_ _1609_ _1610_ _1611_ _1612_ VPWR VGND sg13g2_nor4_1
X_3875_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\] net574 _1544_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_934 VPWR VGND sg13g2_decap_8
XFILLER_32_783 VPWR VGND sg13g2_decap_4
X_2826_ _0759_ _0720_ _0757_ VPWR VGND sg13g2_nand2_2
XFILLER_31_293 VPWR VGND sg13g2_fill_1
X_2757_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[3\] net756 _0741_ _0545_
+ VPWR VGND sg13g2_mux2_1
X_2688_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\] _0723_ _0596_
+ VPWR VGND sg13g2_mux2_1
X_4427_ _2064_ _2068_ _0611_ VPWR VGND sg13g2_nor2_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_24_1018 VPWR VGND sg13g2_decap_8
X_4358_ _2004_ _1999_ _2003_ VPWR VGND sg13g2_xnor2_1
X_3309_ _0999_ videogen.fancy_shader.n646\[4\] videogen.fancy_shader.video_x\[4\]
+ VPWR VGND sg13g2_xnor2_1
X_4289_ _1951_ _1913_ _1923_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_308 VPWR VGND sg13g2_decap_4
XFILLER_39_382 VPWR VGND sg13g2_decap_8
XFILLER_27_533 VPWR VGND sg13g2_decap_8
XFILLER_42_525 VPWR VGND sg13g2_fill_1
XFILLER_42_514 VPWR VGND sg13g2_fill_2
XFILLER_14_205 VPWR VGND sg13g2_decap_4
XFILLER_14_249 VPWR VGND sg13g2_fill_1
XFILLER_11_945 VPWR VGND sg13g2_decap_8
XFILLER_7_927 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_fill_2
XFILLER_6_437 VPWR VGND sg13g2_decap_4
XFILLER_2_643 VPWR VGND sg13g2_decap_8
XFILLER_1_186 VPWR VGND sg13g2_fill_2
XFILLER_49_157 VPWR VGND sg13g2_decap_8
XFILLER_37_319 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_fill_1
XFILLER_46_853 VPWR VGND sg13g2_decap_8
XFILLER_14_761 VPWR VGND sg13g2_fill_2
X_3660_ _1325_ _1326_ _1327_ _1328_ _1329_ VPWR VGND sg13g2_nor4_1
X_2611_ VPWR _0667_ hsync VGND sg13g2_inv_1
X_3591_ _1250_ VPWR _1260_ VGND _1253_ _1258_ sg13g2_o21ai_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_5_481 VPWR VGND sg13g2_fill_1
X_4212_ _1073_ _1870_ _1874_ VPWR VGND sg13g2_nor2_1
X_5192_ net179 VGND VPWR _0616_ blue_tmds_par\[7\] net637 sg13g2_dfrbpq_1
X_5009__226 VPWR VGND net226 sg13g2_tiehi
X_4143_ VPWR _1805_ _1804_ VGND sg13g2_inv_1
X_4074_ _1732_ _1729_ _1739_ VPWR VGND sg13g2_xor2_1
XFILLER_37_820 VPWR VGND sg13g2_fill_1
X_3025_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ _0819_ _0820_ _0821_ VPWR VGND sg13g2_nor4_1
XFILLER_36_363 VPWR VGND sg13g2_decap_8
XFILLER_37_897 VPWR VGND sg13g2_decap_8
X_4976_ net294 VGND VPWR _0404_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[3\]
+ _0061_ sg13g2_dfrbpq_1
X_3927_ VGND VPWR net797 _1298_ _1596_ _1595_ sg13g2_a21oi_1
X_3858_ _1526_ VPWR _1527_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\]
+ net556 sg13g2_o21ai_1
X_3789_ net617 _1452_ _1457_ _1458_ VPWR VGND sg13g2_nor3_1
X_2809_ _0754_ _0699_ _0716_ VPWR VGND sg13g2_nand2_2
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_352 VPWR VGND sg13g2_fill_2
XFILLER_42_300 VPWR VGND sg13g2_decap_4
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_15_558 VPWR VGND sg13g2_decap_4
XFILLER_11_775 VPWR VGND sg13g2_fill_1
X_4856__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_7_768 VPWR VGND sg13g2_fill_2
XFILLER_3_941 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
X_4830_ net650 net702 _0258_ VPWR VGND sg13g2_nor2_1
XFILLER_33_322 VPWR VGND sg13g2_fill_1
XFILLER_33_333 VPWR VGND sg13g2_decap_8
XFILLER_14_591 VPWR VGND sg13g2_decap_4
X_4761_ net668 net719 _0191_ VPWR VGND sg13g2_nor2_1
X_3712_ _1377_ _1378_ _1379_ _1380_ _1381_ VPWR VGND sg13g2_nor4_1
X_4692_ net680 net730 _0122_ VPWR VGND sg13g2_nor2_1
X_3643_ net625 _1306_ _1311_ _1312_ VPWR VGND sg13g2_nor3_1
X_3574_ _1232_ VPWR _1243_ VGND _1236_ _1242_ sg13g2_o21ai_1
X_5244_ net805 VGND VPWR serialize.n427\[5\] serialize.n411\[3\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
Xhold29 serialize.n429\[3\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold18 serialize.n414\[0\] VPWR VGND net423 sg13g2_dlygate4sd3_1
X_5175_ net74 VGND VPWR _0599_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\]
+ _0247_ sg13g2_dfrbpq_1
X_4126_ _1592_ VPWR _1791_ VGND _1398_ _1591_ sg13g2_o21ai_1
XFILLER_37_650 VPWR VGND sg13g2_fill_1
X_4057_ _1722_ _1135_ _1137_ _1720_ VPWR VGND sg13g2_and3_2
X_3008_ _0805_ net629 _0680_ VPWR VGND sg13g2_nand2_1
XFILLER_24_388 VPWR VGND sg13g2_decap_4
X_4959_ net325 VGND VPWR _0387_ red_tmds_par\[8\] net636 sg13g2_dfrbpq_1
XFILLER_10_20 VPWR VGND sg13g2_decap_8
XFILLER_10_53 VPWR VGND sg13g2_fill_1
XFILLER_3_259 VPWR VGND sg13g2_decap_8
XFILLER_0_922 VPWR VGND sg13g2_decap_8
XFILLER_0_999 VPWR VGND sg13g2_decap_8
XFILLER_19_149 VPWR VGND sg13g2_decap_8
XFILLER_28_650 VPWR VGND sg13g2_fill_2
XFILLER_34_119 VPWR VGND sg13g2_decap_4
XFILLER_42_130 VPWR VGND sg13g2_fill_1
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_815 VPWR VGND sg13g2_decap_4
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_15_399 VPWR VGND sg13g2_decap_8
XFILLER_7_510 VPWR VGND sg13g2_decap_4
XFILLER_11_561 VPWR VGND sg13g2_decap_8
XFILLER_7_576 VPWR VGND sg13g2_fill_1
XFILLER_7_565 VPWR VGND sg13g2_decap_8
XFILLER_3_771 VPWR VGND sg13g2_fill_2
X_3290_ net798 VPWR _0983_ VGND videogen.fancy_shader.n646\[1\] _0981_ sg13g2_o21ai_1
XFILLER_25_4 VPWR VGND sg13g2_decap_4
XFILLER_18_160 VPWR VGND sg13g2_decap_8
XFILLER_25_119 VPWR VGND sg13g2_decap_8
XFILLER_46_480 VPWR VGND sg13g2_decap_8
XFILLER_33_141 VPWR VGND sg13g2_fill_1
XFILLER_33_163 VPWR VGND sg13g2_fill_2
X_4813_ net689 net743 _0243_ VPWR VGND sg13g2_nor2_1
XFILLER_22_848 VPWR VGND sg13g2_decap_8
X_4744_ net674 net725 _0174_ VPWR VGND sg13g2_nor2_1
XFILLER_30_892 VPWR VGND sg13g2_fill_1
X_4675_ net684 net737 _0105_ VPWR VGND sg13g2_nor2_1
X_3626_ _1295_ _1238_ _1245_ VPWR VGND sg13g2_nand2_1
X_3557_ VGND VPWR _1226_ _1225_ _1224_ sg13g2_or2_1
X_5227_ net804 VGND VPWR serialize.n429\[1\] serialize.n458 clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3488_ _1150_ _1151_ _1152_ _1153_ _1157_ VPWR VGND sg13g2_and4_1
XFILLER_0_229 VPWR VGND sg13g2_fill_1
X_5158_ net266 VGND VPWR _0582_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\]
+ _0230_ sg13g2_dfrbpq_1
XFILLER_29_414 VPWR VGND sg13g2_decap_4
XFILLER_45_907 VPWR VGND sg13g2_decap_8
X_4109_ _1745_ VPWR _1774_ VGND _1705_ _1753_ sg13g2_o21ai_1
X_5089_ net355 VGND VPWR _0513_ tmds_red.dc_balancing_reg\[4\] net644 sg13g2_dfrbpq_2
XFILLER_44_439 VPWR VGND sg13g2_fill_1
XFILLER_44_428 VPWR VGND sg13g2_decap_4
XFILLER_37_491 VPWR VGND sg13g2_decap_8
XFILLER_12_314 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_fill_2
XFILLER_13_848 VPWR VGND sg13g2_decap_8
XFILLER_9_819 VPWR VGND sg13g2_fill_2
XFILLER_20_380 VPWR VGND sg13g2_fill_1
XFILLER_21_30 VPWR VGND sg13g2_decap_8
X_5150__351 VPWR VGND net351 sg13g2_tiehi
XFILLER_21_96 VPWR VGND sg13g2_decap_8
XFILLER_0_796 VPWR VGND sg13g2_decap_8
XFILLER_47_288 VPWR VGND sg13g2_fill_2
XFILLER_16_653 VPWR VGND sg13g2_decap_4
XFILLER_16_664 VPWR VGND sg13g2_fill_1
X_5040__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_43_472 VPWR VGND sg13g2_fill_2
X_2790_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\] net758 _0750_ _0521_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_852 VPWR VGND sg13g2_fill_1
X_4460_ _2094_ _2079_ _2095_ VPWR VGND sg13g2_xor2_1
X_3411_ _1080_ _1079_ _1078_ VPWR VGND sg13g2_nand2b_1
X_4391_ _2019_ _2035_ _2036_ VPWR VGND sg13g2_and2_1
X_3342_ _1028_ videogen.fancy_shader.n646\[8\] _1026_ VPWR VGND sg13g2_nand2_1
X_3273_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] _0971_ _0973_ VPWR
+ VGND sg13g2_and2_1
X_5012_ net220 VGND VPWR _0440_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\]
+ _0097_ sg13g2_dfrbpq_1
XFILLER_27_907 VPWR VGND sg13g2_decap_8
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_42_29 VPWR VGND sg13g2_decap_8
X_2988_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\] _0800_ _0290_
+ VPWR VGND sg13g2_mux2_1
X_4727_ net650 net703 _0157_ VPWR VGND sg13g2_nor2_1
X_4658_ net667 net720 _0088_ VPWR VGND sg13g2_nor2_1
X_3609_ _1277_ _1263_ _1278_ VPWR VGND sg13g2_xor2_1
X_4589_ net685 net737 _0019_ VPWR VGND sg13g2_nor2_1
XFILLER_27_1005 VPWR VGND sg13g2_decap_8
XFILLER_26_951 VPWR VGND sg13g2_decap_8
XFILLER_25_450 VPWR VGND sg13g2_decap_8
XFILLER_25_461 VPWR VGND sg13g2_decap_8
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_16_85 VPWR VGND sg13g2_fill_2
XFILLER_5_833 VPWR VGND sg13g2_decap_8
X_4974__298 VPWR VGND net298 sg13g2_tiehi
XFILLER_5_888 VPWR VGND sg13g2_decap_8
XFILLER_4_376 VPWR VGND sg13g2_fill_2
XFILLER_4_387 VPWR VGND sg13g2_fill_1
XFILLER_0_571 VPWR VGND sg13g2_decap_8
XFILLER_48_531 VPWR VGND sg13g2_decap_8
XFILLER_36_748 VPWR VGND sg13g2_fill_1
XFILLER_17_940 VPWR VGND sg13g2_decap_8
X_3960_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\] net584 _1628_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_16_450 VPWR VGND sg13g2_fill_2
X_2911_ _0780_ _0716_ _0771_ VPWR VGND sg13g2_nand2_2
XFILLER_32_943 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
X_3891_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\] net550 _1560_ VPWR
+ VGND sg13g2_nor2_1
X_2842_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\] _0762_ _0472_
+ VPWR VGND sg13g2_mux2_1
X_2773_ net790 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\] _0746_ _0534_
+ VPWR VGND sg13g2_mux2_1
X_4512_ _2142_ tmds_blue.dc_balancing_reg\[2\] _2140_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_693 VPWR VGND sg13g2_decap_8
X_4443_ _2079_ net600 _2077_ _2078_ VPWR VGND sg13g2_and3_2
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
X_4374_ _0910_ _2018_ _2019_ _2020_ VPWR VGND sg13g2_nor3_1
Xfanout628 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[0\] net628 VPWR VGND
+ sg13g2_buf_8
X_3325_ VGND VPWR _1002_ _1006_ _1015_ _1001_ sg13g2_a21oi_1
Xfanout639 net640 net639 VPWR VGND sg13g2_buf_8
Xfanout617 videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\] net617 VPWR VGND
+ sg13g2_buf_8
X_3256_ _0809_ _0961_ _0326_ VPWR VGND sg13g2_nor2_1
XFILLER_39_531 VPWR VGND sg13g2_decap_8
XFILLER_39_564 VPWR VGND sg13g2_fill_2
X_3187_ VGND VPWR tmds_red.n100 _0914_ _0274_ _0915_ sg13g2_a21oi_1
XFILLER_26_214 VPWR VGND sg13g2_decap_4
XFILLER_26_225 VPWR VGND sg13g2_decap_8
XFILLER_27_737 VPWR VGND sg13g2_decap_8
XFILLER_27_748 VPWR VGND sg13g2_fill_1
XFILLER_42_707 VPWR VGND sg13g2_fill_1
XFILLER_14_409 VPWR VGND sg13g2_decap_4
XFILLER_22_420 VPWR VGND sg13g2_fill_2
XFILLER_23_965 VPWR VGND sg13g2_decap_8
X_5019__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_2_803 VPWR VGND sg13g2_decap_8
XFILLER_1_313 VPWR VGND sg13g2_fill_2
XFILLER_40_1013 VPWR VGND sg13g2_decap_8
XFILLER_17_203 VPWR VGND sg13g2_decap_4
XFILLER_18_748 VPWR VGND sg13g2_fill_1
XFILLER_18_759 VPWR VGND sg13g2_fill_1
XFILLER_14_910 VPWR VGND sg13g2_decap_8
XFILLER_43_50 VPWR VGND sg13g2_decap_4
XFILLER_9_402 VPWR VGND sg13g2_decap_8
XFILLER_9_435 VPWR VGND sg13g2_fill_2
XFILLER_13_453 VPWR VGND sg13g2_decap_8
XFILLER_14_987 VPWR VGND sg13g2_decap_8
XFILLER_5_630 VPWR VGND sg13g2_fill_1
X_3110_ red_tmds_par\[8\] net695 serialize.n427\[8\] VPWR VGND sg13g2_and2_1
X_4866__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_0_390 VPWR VGND sg13g2_decap_8
X_4090_ _1755_ _1065_ _0990_ VPWR VGND sg13g2_nand2b_1
X_3041_ _0683_ _0694_ _0828_ VPWR VGND sg13g2_nor2_1
XFILLER_48_394 VPWR VGND sg13g2_decap_8
X_5120__209 VPWR VGND net209 sg13g2_tiehi
X_4992_ net259 VGND VPWR _0420_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[3\]
+ _0077_ sg13g2_dfrbpq_1
XFILLER_17_792 VPWR VGND sg13g2_decap_8
XFILLER_16_291 VPWR VGND sg13g2_fill_1
XFILLER_32_740 VPWR VGND sg13g2_decap_8
X_3943_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\] net558 _1611_ VPWR
+ VGND sg13g2_nor2_1
X_3874_ net620 VPWR _1543_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[3\]
+ net584 sg13g2_o21ai_1
XFILLER_20_913 VPWR VGND sg13g2_decap_8
X_2825_ _0758_ net545 _0743_ VPWR VGND sg13g2_nand2_2
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_2756_ _0707_ _0733_ _0741_ VPWR VGND sg13g2_nor2_2
X_2687_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\] _0723_ _0597_
+ VPWR VGND sg13g2_mux2_1
X_4426_ tmds_blue.dc_balancing_reg\[4\] _2067_ _2068_ VPWR VGND sg13g2_nor2_2
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4357_ VPWR _2003_ _2002_ VGND sg13g2_inv_1
X_3308_ _0998_ videogen.fancy_shader.n646\[4\] videogen.fancy_shader.video_x\[4\]
+ VPWR VGND sg13g2_nand2_1
X_4288_ _1942_ _1943_ _1925_ _1950_ VPWR VGND _1945_ sg13g2_nand4_1
X_3239_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0948_ _0950_ VPWR VGND
+ sg13g2_and2_1
XFILLER_42_504 VPWR VGND sg13g2_decap_4
XFILLER_27_578 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_decap_8
XFILLER_42_559 VPWR VGND sg13g2_decap_8
XFILLER_42_548 VPWR VGND sg13g2_fill_1
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_7_906 VPWR VGND sg13g2_decap_8
XFILLER_13_75 VPWR VGND sg13g2_decap_8
XFILLER_10_489 VPWR VGND sg13g2_fill_1
X_4905__40 VPWR VGND net40 sg13g2_tiehi
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_49_114 VPWR VGND sg13g2_decap_8
XFILLER_2_677 VPWR VGND sg13g2_decap_8
XFILLER_18_501 VPWR VGND sg13g2_decap_8
XFILLER_18_512 VPWR VGND sg13g2_fill_1
XFILLER_18_534 VPWR VGND sg13g2_fill_1
XFILLER_13_283 VPWR VGND sg13g2_fill_1
X_3590_ VGND VPWR _1259_ _1258_ _1253_ sg13g2_or2_1
X_2610_ VPWR _0666_ tmds_red.dc_balancing_reg\[3\] VGND sg13g2_inv_1
XFILLER_5_471 VPWR VGND sg13g2_decap_4
X_4211_ VPWR _1873_ _1872_ VGND sg13g2_inv_1
X_5191_ net187 VGND VPWR _0615_ blue_tmds_par\[6\] net637 sg13g2_dfrbpq_1
X_4142_ _1804_ _1718_ _1802_ VPWR VGND sg13g2_xnor2_1
X_4073_ _1738_ _1735_ _1737_ _1732_ _1730_ VPWR VGND sg13g2_a22oi_1
X_3024_ VGND VPWR _0820_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\]
+ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\] sg13g2_or2_1
XFILLER_24_515 VPWR VGND sg13g2_fill_1
X_4975_ net296 VGND VPWR _0403_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\]
+ _0060_ sg13g2_dfrbpq_1
X_3926_ _1496_ _1594_ _1595_ VPWR VGND sg13g2_nor2_1
X_3857_ _1526_ net583 _0633_ net594 _0632_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
X_3788_ net625 _1453_ _1454_ _1456_ _1457_ VPWR VGND sg13g2_nor4_1
X_2808_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\] net784 _0753_ _0497_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_787 VPWR VGND sg13g2_decap_8
X_2739_ net794 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\] _0736_ _0558_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
X_4409_ VGND VPWR _2030_ _2051_ _2053_ _2052_ sg13g2_a21oi_1
XFILLER_28_810 VPWR VGND sg13g2_decap_4
XFILLER_39_180 VPWR VGND sg13g2_decap_8
XFILLER_27_342 VPWR VGND sg13g2_fill_2
XFILLER_30_518 VPWR VGND sg13g2_fill_2
XFILLER_11_721 VPWR VGND sg13g2_fill_1
XFILLER_7_714 VPWR VGND sg13g2_decap_8
XFILLER_6_202 VPWR VGND sg13g2_fill_2
XFILLER_40_40 VPWR VGND sg13g2_fill_2
XFILLER_6_268 VPWR VGND sg13g2_fill_1
XFILLER_3_920 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_4
XFILLER_3_997 VPWR VGND sg13g2_decap_8
XFILLER_38_618 VPWR VGND sg13g2_fill_1
XFILLER_19_821 VPWR VGND sg13g2_fill_1
XFILLER_19_876 VPWR VGND sg13g2_decap_4
XFILLER_46_684 VPWR VGND sg13g2_fill_2
X_4760_ net668 net723 _0190_ VPWR VGND sg13g2_nor2_1
X_3711_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\] net578 _1380_ VPWR
+ VGND sg13g2_nor2_1
X_4691_ net675 net727 _0121_ VPWR VGND sg13g2_nor2_1
X_3642_ _1307_ _1308_ _1309_ _1310_ _1311_ VPWR VGND sg13g2_nor4_1
X_3573_ _1242_ _1238_ _1240_ _1241_ VPWR VGND sg13g2_and3_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_5243_ net802 VGND VPWR serialize.n427\[4\] serialize.n411\[2\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
Xhold19 serialize.n411\[3\] VPWR VGND net424 sg13g2_dlygate4sd3_1
X_5174_ net100 VGND VPWR _0598_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\]
+ _0246_ sg13g2_dfrbpq_1
X_4125_ _1297_ VPWR _1790_ VGND _1783_ _1789_ sg13g2_o21ai_1
X_5206__250 VPWR VGND net250 sg13g2_tiehi
X_4056_ VGND VPWR _1720_ _1721_ _1137_ _1135_ sg13g2_a21oi_2
X_3007_ net629 _0680_ _0804_ VPWR VGND sg13g2_and2_1
XFILLER_24_301 VPWR VGND sg13g2_fill_1
XFILLER_25_835 VPWR VGND sg13g2_decap_8
X_5073__31 VPWR VGND net31 sg13g2_tiehi
XFILLER_25_879 VPWR VGND sg13g2_decap_8
X_4958_ net326 VGND VPWR _0386_ red_tmds_par\[6\] net641 sg13g2_dfrbpq_1
XFILLER_20_551 VPWR VGND sg13g2_decap_8
X_4889_ net71 VGND VPWR _0317_ tmds_blue.vsync net636 sg13g2_dfrbpq_1
X_3909_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\] net580 _1578_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_10_76 VPWR VGND sg13g2_fill_2
XFILLER_0_901 VPWR VGND sg13g2_decap_8
X_4887__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_27_150 VPWR VGND sg13g2_decap_8
XFILLER_37_1007 VPWR VGND sg13g2_decap_8
XFILLER_16_868 VPWR VGND sg13g2_fill_2
XFILLER_27_194 VPWR VGND sg13g2_fill_2
XFILLER_7_522 VPWR VGND sg13g2_decap_8
XFILLER_7_544 VPWR VGND sg13g2_decap_8
XFILLER_3_794 VPWR VGND sg13g2_decap_8
X_4984__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_38_426 VPWR VGND sg13g2_decap_8
XFILLER_38_459 VPWR VGND sg13g2_fill_2
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
XFILLER_21_337 VPWR VGND sg13g2_decap_8
X_4812_ net689 net739 _0242_ VPWR VGND sg13g2_nor2_1
XFILLER_33_175 VPWR VGND sg13g2_fill_2
XFILLER_34_698 VPWR VGND sg13g2_decap_8
X_4743_ net656 net708 _0173_ VPWR VGND sg13g2_nor2_1
X_4674_ net686 net738 _0104_ VPWR VGND sg13g2_nor2_1
X_3625_ _1287_ _1293_ _1294_ VPWR VGND sg13g2_nor2b_1
X_3556_ _1225_ _1189_ _1208_ _1223_ VPWR VGND sg13g2_and3_1
X_5226_ net804 VGND VPWR serialize.n429\[0\] serialize.n456 clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3487_ _1156_ _1152_ _1153_ _1151_ _1150_ VPWR VGND sg13g2_a22oi_1
X_5157_ net273 VGND VPWR _0581_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\]
+ _0229_ sg13g2_dfrbpq_1
X_4108_ VPWR VGND _1765_ _1754_ _1763_ _1755_ _1773_ _1756_ sg13g2_a221oi_1
X_5088_ net357 VGND VPWR _0512_ tmds_red.dc_balancing_reg\[3\] net644 sg13g2_dfrbpq_1
XFILLER_38_993 VPWR VGND sg13g2_decap_8
X_4039_ _1704_ _0995_ _1195_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_602 VPWR VGND sg13g2_fill_1
XFILLER_24_131 VPWR VGND sg13g2_decap_8
XFILLER_25_654 VPWR VGND sg13g2_fill_1
XFILLER_40_635 VPWR VGND sg13g2_fill_1
XFILLER_24_164 VPWR VGND sg13g2_decap_8
XFILLER_24_175 VPWR VGND sg13g2_fill_1
XFILLER_12_359 VPWR VGND sg13g2_decap_4
XFILLER_20_370 VPWR VGND sg13g2_fill_2
XFILLER_4_514 VPWR VGND sg13g2_fill_2
XFILLER_4_503 VPWR VGND sg13g2_decap_8
XFILLER_43_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
XFILLER_47_256 VPWR VGND sg13g2_decap_4
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_16_621 VPWR VGND sg13g2_fill_2
XFILLER_44_985 VPWR VGND sg13g2_decap_8
XFILLER_43_440 VPWR VGND sg13g2_fill_2
XFILLER_15_142 VPWR VGND sg13g2_decap_8
XFILLER_31_602 VPWR VGND sg13g2_fill_2
XFILLER_15_186 VPWR VGND sg13g2_decap_8
XFILLER_30_101 VPWR VGND sg13g2_fill_2
XFILLER_30_134 VPWR VGND sg13g2_decap_8
X_5116__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_7_352 VPWR VGND sg13g2_decap_4
X_3410_ _1079_ videogen.fancy_shader.n646\[5\] videogen.fancy_shader.video_x\[5\]
+ VPWR VGND sg13g2_nand2_1
X_4390_ _2035_ _2031_ _2033_ VPWR VGND sg13g2_xnor2_1
X_3341_ VGND VPWR _1027_ _1026_ net609 sg13g2_or2_1
XFILLER_3_591 VPWR VGND sg13g2_decap_4
X_3272_ VGND VPWR _0938_ _0971_ _0972_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[2\]
+ sg13g2_a21oi_1
X_5011_ net222 VGND VPWR _0439_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\]
+ _0096_ sg13g2_dfrbpq_1
XFILLER_39_757 VPWR VGND sg13g2_decap_4
XFILLER_38_278 VPWR VGND sg13g2_decap_8
XFILLER_26_407 VPWR VGND sg13g2_decap_4
XFILLER_26_429 VPWR VGND sg13g2_fill_1
XFILLER_34_440 VPWR VGND sg13g2_decap_4
X_2987_ _0800_ _0722_ _0771_ VPWR VGND sg13g2_nand2_2
XFILLER_21_156 VPWR VGND sg13g2_decap_8
X_4726_ net654 net705 _0156_ VPWR VGND sg13g2_nor2_1
X_4657_ net669 net722 _0087_ VPWR VGND sg13g2_nor2_1
X_3608_ VGND VPWR _1268_ _1273_ _1277_ _1266_ sg13g2_a21oi_1
X_4588_ net685 net737 _0018_ VPWR VGND sg13g2_nor2_1
X_3539_ _1206_ _1201_ _1195_ _1208_ VPWR VGND sg13g2_a21o_1
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
X_5209_ net803 VGND VPWR serialize.n428\[1\] serialize.n455 clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_18_919 VPWR VGND sg13g2_decap_8
XFILLER_44_226 VPWR VGND sg13g2_fill_1
XFILLER_26_930 VPWR VGND sg13g2_decap_8
XFILLER_41_922 VPWR VGND sg13g2_fill_2
XFILLER_41_911 VPWR VGND sg13g2_decap_4
XFILLER_13_624 VPWR VGND sg13g2_fill_2
XFILLER_16_97 VPWR VGND sg13g2_decap_8
XFILLER_40_465 VPWR VGND sg13g2_decap_8
XFILLER_12_189 VPWR VGND sg13g2_decap_4
XFILLER_10_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_867 VPWR VGND sg13g2_decap_8
XFILLER_0_550 VPWR VGND sg13g2_decap_8
XFILLER_36_716 VPWR VGND sg13g2_fill_1
XFILLER_35_204 VPWR VGND sg13g2_fill_2
X_2910_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\] net788 _0779_ _0421_
+ VPWR VGND sg13g2_mux2_1
XFILLER_44_793 VPWR VGND sg13g2_fill_2
XFILLER_17_996 VPWR VGND sg13g2_decap_8
XFILLER_32_922 VPWR VGND sg13g2_decap_8
X_3890_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\] net574 _1559_ VPWR
+ VGND sg13g2_nor2_1
X_2841_ _0762_ _0711_ _0757_ VPWR VGND sg13g2_nand2_2
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_2772_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\] _0746_ _0535_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_672 VPWR VGND sg13g2_fill_2
XFILLER_8_661 VPWR VGND sg13g2_decap_8
X_4511_ _2141_ _2140_ tmds_blue.dc_balancing_reg\[2\] VPWR VGND sg13g2_nand2b_1
X_4442_ _2078_ net599 _0652_ VPWR VGND sg13g2_nand2_1
X_4373_ _2012_ _2017_ _2019_ VPWR VGND sg13g2_nor2_1
Xfanout629 videogen.fancy_shader.video_x\[7\] net629 VPWR VGND sg13g2_buf_8
X_3324_ _1014_ videogen.fancy_shader.n646\[3\] videogen.fancy_shader.video_x\[3\]
+ VPWR VGND sg13g2_xnor2_1
Xfanout618 net620 net618 VPWR VGND sg13g2_buf_8
Xfanout607 display_enable net607 VPWR VGND sg13g2_buf_8
X_3255_ _0961_ net623 _0959_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_204 VPWR VGND sg13g2_fill_1
X_3186_ _0852_ VPWR _0915_ VGND tmds_red.n100 _0914_ sg13g2_o21ai_1
XFILLER_22_410 VPWR VGND sg13g2_decap_4
XFILLER_35_771 VPWR VGND sg13g2_decap_8
XFILLER_23_944 VPWR VGND sg13g2_decap_8
X_4709_ net680 net732 _0139_ VPWR VGND sg13g2_nor2_1
XFILLER_2_859 VPWR VGND sg13g2_decap_8
XFILLER_18_705 VPWR VGND sg13g2_decap_8
X_5106__268 VPWR VGND net268 sg13g2_tiehi
XFILLER_27_74 VPWR VGND sg13g2_fill_2
XFILLER_26_760 VPWR VGND sg13g2_fill_2
XFILLER_26_771 VPWR VGND sg13g2_decap_8
XFILLER_14_966 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_fill_1
XFILLER_5_686 VPWR VGND sg13g2_fill_1
XFILLER_4_196 VPWR VGND sg13g2_fill_1
XFILLER_4_45 VPWR VGND sg13g2_decap_8
XFILLER_48_362 VPWR VGND sg13g2_fill_1
X_3040_ VGND VPWR net595 net13 _0695_ net549 sg13g2_a21oi_2
XFILLER_49_896 VPWR VGND sg13g2_decap_8
XFILLER_36_535 VPWR VGND sg13g2_fill_1
XFILLER_36_579 VPWR VGND sg13g2_decap_8
X_4991_ net265 VGND VPWR _0419_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\]
+ _0076_ sg13g2_dfrbpq_1
XFILLER_17_760 VPWR VGND sg13g2_fill_1
XFILLER_23_218 VPWR VGND sg13g2_decap_8
X_3942_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\] net568 _1610_ VPWR
+ VGND sg13g2_nor2_1
X_3873_ _1519_ _1541_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1542_
+ VPWR VGND sg13g2_nand3_1
X_2824_ net545 _0743_ _0757_ VPWR VGND sg13g2_and2_1
XFILLER_20_969 VPWR VGND sg13g2_decap_8
X_2755_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\] net786 _0740_ _0546_
+ VPWR VGND sg13g2_mux2_1
X_2686_ _0723_ _0722_ VPWR VGND _0719_ sg13g2_nand2b_2
X_4425_ net605 VPWR _2067_ VGND _2056_ _2066_ sg13g2_o21ai_1
X_4356_ VGND VPWR _0665_ _0869_ _2002_ _2001_ sg13g2_a21oi_1
X_3307_ net750 _0997_ _0349_ VPWR VGND sg13g2_nor2_1
X_4287_ _1949_ _1942_ _1943_ VPWR VGND sg13g2_nand2_1
X_3238_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\] _0948_ _0949_ VPWR VGND
+ sg13g2_nor2_1
X_3169_ _0897_ _0896_ _0898_ VPWR VGND sg13g2_xor2_1
XFILLER_15_708 VPWR VGND sg13g2_decap_4
XFILLER_42_516 VPWR VGND sg13g2_fill_1
XFILLER_11_903 VPWR VGND sg13g2_decap_8
XFILLER_23_796 VPWR VGND sg13g2_fill_2
XFILLER_38_51 VPWR VGND sg13g2_fill_1
XFILLER_18_546 VPWR VGND sg13g2_decap_8
XFILLER_46_888 VPWR VGND sg13g2_decap_8
XFILLER_45_398 VPWR VGND sg13g2_decap_4
XFILLER_33_538 VPWR VGND sg13g2_fill_2
XFILLER_41_571 VPWR VGND sg13g2_fill_1
XFILLER_6_984 VPWR VGND sg13g2_decap_8
X_4210_ _1872_ _1838_ _1871_ VPWR VGND sg13g2_xnor2_1
X_5190_ net195 VGND VPWR _0614_ blue_tmds_par\[5\] net638 sg13g2_dfrbpq_1
X_4141_ _1082_ _1142_ _1018_ _1803_ VPWR VGND sg13g2_nand3_1
X_4072_ _1729_ _1732_ _1728_ _1737_ VPWR VGND sg13g2_nand3_1
X_3023_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\]
+ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] _0819_ VPWR VGND sg13g2_nand3_1
XFILLER_24_527 VPWR VGND sg13g2_decap_4
X_4974_ net298 VGND VPWR _0402_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\]
+ _0059_ sg13g2_dfrbpq_1
XFILLER_17_590 VPWR VGND sg13g2_fill_1
X_3925_ _1594_ net797 _1593_ VPWR VGND sg13g2_nand2_1
XFILLER_32_582 VPWR VGND sg13g2_fill_2
X_3856_ net616 VPWR _1525_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\]
+ net570 sg13g2_o21ai_1
X_3787_ _1455_ VPWR _1456_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\]
+ net558 sg13g2_o21ai_1
X_2807_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\] net773 _0753_ _0498_
+ VPWR VGND sg13g2_mux2_1
X_2738_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\] _0736_ _0559_
+ VPWR VGND sg13g2_mux2_1
X_2669_ VGND VPWR _0714_ _0698_ net545 sg13g2_or2_1
X_4408_ _0910_ VPWR _2052_ VGND _2030_ _2051_ sg13g2_o21ai_1
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
X_4339_ net747 _1991_ _0388_ VPWR VGND sg13g2_nor2_1
XFILLER_28_855 VPWR VGND sg13g2_decap_4
XFILLER_27_387 VPWR VGND sg13g2_fill_2
XFILLER_42_368 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_24_64 VPWR VGND sg13g2_decap_8
XFILLER_10_232 VPWR VGND sg13g2_fill_2
XFILLER_24_86 VPWR VGND sg13g2_decap_8
XFILLER_6_225 VPWR VGND sg13g2_decap_8
XFILLER_2_420 VPWR VGND sg13g2_decap_8
XFILLER_3_976 VPWR VGND sg13g2_decap_8
Xfanout790 net793 net790 VPWR VGND sg13g2_buf_8
XFILLER_19_855 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_fill_2
XFILLER_45_173 VPWR VGND sg13g2_fill_2
XFILLER_34_847 VPWR VGND sg13g2_decap_8
X_3710_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\] net567 _1379_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_14_1008 VPWR VGND sg13g2_decap_8
X_4690_ net675 net727 _0120_ VPWR VGND sg13g2_nor2_1
X_3641_ videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\] net591 _1310_ VPWR
+ VGND sg13g2_nor2_1
X_4919__384 VPWR VGND net384 sg13g2_tiehi
X_3572_ _1213_ VPWR _1241_ VGND _1219_ _1239_ sg13g2_o21ai_1
XFILLER_5_280 VPWR VGND sg13g2_fill_2
X_5089__355 VPWR VGND net355 sg13g2_tiehi
X_5242_ net802 VGND VPWR serialize.n427\[3\] serialize.n411\[1\] clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_5173_ net116 VGND VPWR _0597_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\]
+ _0245_ sg13g2_dfrbpq_1
X_4124_ _1785_ _1786_ _1784_ _1789_ VPWR VGND _1788_ sg13g2_nand4_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_2
XFILLER_49_490 VPWR VGND sg13g2_decap_8
XFILLER_37_641 VPWR VGND sg13g2_decap_8
X_4055_ _1163_ _1710_ _1720_ VPWR VGND sg13g2_and2_1
X_3006_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\] _0803_ _0267_
+ VPWR VGND sg13g2_mux2_1
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_24_335 VPWR VGND sg13g2_decap_8
XFILLER_25_858 VPWR VGND sg13g2_decap_8
X_4957_ net327 VGND VPWR _0385_ red_tmds_par\[4\] net641 sg13g2_dfrbpq_1
X_4888_ net73 VGND VPWR _0316_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\]
+ _0037_ sg13g2_dfrbpq_1
X_3908_ net625 VPWR _1577_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\]
+ net590 sg13g2_o21ai_1
X_3839_ net598 VPWR _1508_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\]
+ net587 sg13g2_o21ai_1
XFILLER_10_44 VPWR VGND sg13g2_fill_1
XFILLER_0_957 VPWR VGND sg13g2_decap_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_4
XFILLER_19_118 VPWR VGND sg13g2_decap_8
XFILLER_19_129 VPWR VGND sg13g2_fill_2
XFILLER_28_652 VPWR VGND sg13g2_fill_1
XFILLER_43_644 VPWR VGND sg13g2_fill_2
XFILLER_42_121 VPWR VGND sg13g2_decap_8
XFILLER_15_313 VPWR VGND sg13g2_fill_2
XFILLER_15_335 VPWR VGND sg13g2_decap_4
XFILLER_3_773 VPWR VGND sg13g2_fill_1
XFILLER_32_7 VPWR VGND sg13g2_fill_1
XFILLER_39_939 VPWR VGND sg13g2_decap_8
XFILLER_38_405 VPWR VGND sg13g2_fill_2
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_18_195 VPWR VGND sg13g2_decap_4
XFILLER_34_633 VPWR VGND sg13g2_decap_8
XFILLER_22_817 VPWR VGND sg13g2_decap_8
X_4811_ net689 net739 _0241_ VPWR VGND sg13g2_nor2_1
XFILLER_15_891 VPWR VGND sg13g2_decap_8
X_5055__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_33_165 VPWR VGND sg13g2_fill_1
X_4742_ net656 net708 _0172_ VPWR VGND sg13g2_nor2_1
X_4673_ net686 net738 _0103_ VPWR VGND sg13g2_nor2_1
X_3624_ _1293_ _1292_ _1285_ _1289_ _1284_ VPWR VGND sg13g2_a22oi_1
X_3555_ VGND VPWR _1208_ _1223_ _1224_ _1189_ sg13g2_a21oi_1
X_3486_ _1143_ _1098_ _1097_ _1155_ VPWR VGND sg13g2_a21o_1
X_5225_ net800 VGND VPWR net694 serialize.n420\[6\] clknet_3_2__leaf_clk_regs sg13g2_dfrbpq_1
X_5156_ net281 VGND VPWR _0580_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\]
+ _0228_ sg13g2_dfrbpq_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_4963__319 VPWR VGND net319 sg13g2_tiehi
X_4107_ _1769_ _1771_ _1772_ VPWR VGND _1768_ sg13g2_nand3b_1
XFILLER_29_438 VPWR VGND sg13g2_fill_2
X_5087_ net359 VGND VPWR _0511_ tmds_red.dc_balancing_reg\[2\] net644 sg13g2_dfrbpq_2
XFILLER_38_972 VPWR VGND sg13g2_decap_8
X_4038_ _1703_ _1060_ _1702_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_644 VPWR VGND sg13g2_fill_1
XFILLER_24_121 VPWR VGND sg13g2_decap_4
XFILLER_25_677 VPWR VGND sg13g2_decap_8
XFILLER_13_839 VPWR VGND sg13g2_fill_1
XFILLER_21_872 VPWR VGND sg13g2_fill_2
XFILLER_21_76 VPWR VGND sg13g2_decap_8
XFILLER_0_754 VPWR VGND sg13g2_decap_8
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_28_471 VPWR VGND sg13g2_decap_8
XFILLER_44_964 VPWR VGND sg13g2_decap_8
XFILLER_43_496 VPWR VGND sg13g2_fill_2
XFILLER_43_485 VPWR VGND sg13g2_fill_2
XFILLER_43_474 VPWR VGND sg13g2_fill_1
XFILLER_31_658 VPWR VGND sg13g2_decap_8
XFILLER_12_861 VPWR VGND sg13g2_fill_2
XFILLER_8_843 VPWR VGND sg13g2_decap_8
XFILLER_7_331 VPWR VGND sg13g2_fill_1
XFILLER_8_898 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_fill_2
XFILLER_7_386 VPWR VGND sg13g2_fill_1
XFILLER_7_89 VPWR VGND sg13g2_decap_8
X_3340_ net745 _1025_ _1026_ _0353_ VPWR VGND sg13g2_nor3_1
X_5010_ net224 VGND VPWR _0438_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\]
+ _0095_ sg13g2_dfrbpq_1
X_3271_ _0967_ _0970_ _0971_ _0331_ VPWR VGND sg13g2_nor3_1
XFILLER_39_714 VPWR VGND sg13g2_decap_8
XFILLER_38_257 VPWR VGND sg13g2_fill_2
XFILLER_19_493 VPWR VGND sg13g2_decap_8
XFILLER_35_931 VPWR VGND sg13g2_decap_8
XFILLER_35_997 VPWR VGND sg13g2_decap_8
X_5093__318 VPWR VGND net318 sg13g2_tiehi
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_21_135 VPWR VGND sg13g2_fill_2
X_2986_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\] _0799_ _0291_
+ VPWR VGND sg13g2_mux2_1
X_4725_ net651 net702 _0155_ VPWR VGND sg13g2_nor2_1
X_4656_ net669 net722 _0086_ VPWR VGND sg13g2_nor2_1
X_3607_ _1066_ _1273_ _1274_ _1276_ VPWR VGND sg13g2_nor3_1
X_4587_ net657 net709 _0017_ VPWR VGND sg13g2_nor2_1
X_3538_ _1207_ _1200_ _1198_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_529 VPWR VGND sg13g2_decap_8
X_3469_ _1138_ _1135_ _1137_ VPWR VGND sg13g2_nand2_1
X_5208_ net803 VGND VPWR serialize.n428\[0\] serialize.n453 clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_235 VPWR VGND sg13g2_decap_8
X_5139_ net86 VGND VPWR _0563_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\]
+ _0211_ sg13g2_dfrbpq_1
XFILLER_29_257 VPWR VGND sg13g2_decap_4
XFILLER_45_739 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_fill_1
XFILLER_38_791 VPWR VGND sg13g2_fill_2
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_16_65 VPWR VGND sg13g2_fill_1
XFILLER_26_986 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_4
XFILLER_40_444 VPWR VGND sg13g2_decap_8
XFILLER_10_1000 VPWR VGND sg13g2_decap_8
XFILLER_4_378 VPWR VGND sg13g2_fill_1
XFILLER_48_577 VPWR VGND sg13g2_fill_2
XFILLER_48_566 VPWR VGND sg13g2_decap_8
XFILLER_17_975 VPWR VGND sg13g2_decap_8
XFILLER_43_260 VPWR VGND sg13g2_fill_2
XFILLER_16_452 VPWR VGND sg13g2_fill_1
X_2840_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\] _0761_ _0473_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_978 VPWR VGND sg13g2_decap_8
XFILLER_8_640 VPWR VGND sg13g2_fill_1
X_2771_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\] _0746_ _0536_
+ VPWR VGND sg13g2_mux2_1
X_4510_ _2138_ _2139_ _2140_ VPWR VGND sg13g2_nor2_2
X_4441_ _2077_ tmds_green.dc_balancing_reg\[1\] net599 VPWR VGND sg13g2_nand2b_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
X_4372_ _2014_ _2017_ _2018_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_890 VPWR VGND sg13g2_decap_8
Xfanout619 net620 net619 VPWR VGND sg13g2_buf_8
X_3323_ _1011_ _1012_ _1013_ VPWR VGND sg13g2_and2_1
Xfanout608 videogen.fancy_shader.video_y\[0\] net608 VPWR VGND sg13g2_buf_8
XFILLER_39_500 VPWR VGND sg13g2_decap_4
X_3254_ _0809_ _0959_ _0960_ _0325_ VPWR VGND sg13g2_nor3_1
X_3185_ _0912_ _0913_ _0914_ VPWR VGND sg13g2_nor2_2
XFILLER_23_923 VPWR VGND sg13g2_decap_8
XFILLER_34_260 VPWR VGND sg13g2_decap_4
XFILLER_22_422 VPWR VGND sg13g2_fill_1
XFILLER_34_282 VPWR VGND sg13g2_fill_1
XFILLER_35_794 VPWR VGND sg13g2_fill_2
XFILLER_10_617 VPWR VGND sg13g2_fill_2
XFILLER_22_477 VPWR VGND sg13g2_fill_1
X_2969_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\] _0794_ _0313_
+ VPWR VGND sg13g2_mux2_1
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
X_4708_ net680 net730 _0138_ VPWR VGND sg13g2_nor2_1
X_4639_ net664 net716 _0069_ VPWR VGND sg13g2_nor2_1
XFILLER_2_838 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_fill_1
XFILLER_45_569 VPWR VGND sg13g2_decap_8
XFILLER_45_558 VPWR VGND sg13g2_decap_8
XFILLER_32_219 VPWR VGND sg13g2_fill_2
XFILLER_14_945 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_fill_2
XFILLER_5_621 VPWR VGND sg13g2_decap_4
XFILLER_1_893 VPWR VGND sg13g2_decap_8
XFILLER_49_875 VPWR VGND sg13g2_decap_8
XFILLER_24_709 VPWR VGND sg13g2_fill_2
X_4990_ net267 VGND VPWR _0418_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\]
+ _0075_ sg13g2_dfrbpq_1
XFILLER_17_783 VPWR VGND sg13g2_fill_1
XFILLER_23_208 VPWR VGND sg13g2_decap_4
XFILLER_44_591 VPWR VGND sg13g2_fill_1
X_3941_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\] net580 _1609_ VPWR
+ VGND sg13g2_nor2_1
X_3872_ _1540_ VPWR _1541_ VGND _1524_ _1528_ sg13g2_o21ai_1
XFILLER_17_1017 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_32_764 VPWR VGND sg13g2_decap_8
X_2823_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\] net789 _0756_ _0485_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_948 VPWR VGND sg13g2_decap_8
XFILLER_31_274 VPWR VGND sg13g2_decap_8
X_2754_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[1\] net775 _0740_ _0547_
+ VPWR VGND sg13g2_mux2_1
X_2685_ net619 net628 net595 _0722_ VGND VPWR _0705_ sg13g2_nor4_2
X_4424_ _2066_ net604 tmds_blue.n193 VPWR VGND sg13g2_xnor2_1
X_4355_ _0869_ _0898_ _2001_ VPWR VGND sg13g2_nor2_1
X_3306_ _0997_ videogen.fancy_shader.n646\[3\] _0996_ VPWR VGND sg13g2_xnor2_1
X_4286_ _1937_ _1947_ _1948_ VPWR VGND sg13g2_nor2_1
XFILLER_39_341 VPWR VGND sg13g2_decap_4
X_3237_ _0943_ _0947_ _0948_ _0320_ VPWR VGND sg13g2_nor3_1
X_4929__364 VPWR VGND net364 sg13g2_tiehi
XFILLER_39_363 VPWR VGND sg13g2_decap_8
X_3168_ VGND VPWR tmds_red.n102 _0885_ _0897_ _0887_ sg13g2_a21oi_1
XFILLER_27_547 VPWR VGND sg13g2_fill_2
X_3099_ net438 green_tmds_par\[7\] net698 serialize.n428\[7\] VPWR VGND sg13g2_mux2_1
X_5179__381 VPWR VGND net381 sg13g2_tiehi
XFILLER_10_425 VPWR VGND sg13g2_fill_1
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_6_407 VPWR VGND sg13g2_fill_2
XFILLER_13_44 VPWR VGND sg13g2_decap_8
XFILLER_13_55 VPWR VGND sg13g2_fill_2
X_5112__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_38_74 VPWR VGND sg13g2_decap_8
XFILLER_46_867 VPWR VGND sg13g2_decap_8
XFILLER_14_720 VPWR VGND sg13g2_fill_2
XFILLER_9_289 VPWR VGND sg13g2_fill_2
XFILLER_6_963 VPWR VGND sg13g2_decap_8
X_4140_ _1802_ _1018_ _1082_ VPWR VGND sg13g2_nand2_2
X_4071_ _1736_ _1729_ _1732_ VPWR VGND sg13g2_nand2_1
XFILLER_23_1021 VPWR VGND sg13g2_decap_8
X_3022_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0807_ _0818_ VPWR
+ VGND sg13g2_and2_1
X_4973_ net300 VGND VPWR _0401_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[0\]
+ _0058_ sg13g2_dfrbpq_1
X_3924_ net1 _1591_ _1593_ VPWR VGND sg13g2_nor2_1
X_3855_ _1520_ _1521_ _1522_ _1523_ _1524_ VPWR VGND sg13g2_nor4_1
XFILLER_20_745 VPWR VGND sg13g2_decap_8
X_3786_ _1455_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
X_2806_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\] net762 _0753_ _0499_
+ VPWR VGND sg13g2_mux2_1
X_2737_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\] _0736_ _0560_
+ VPWR VGND sg13g2_mux2_1
X_2668_ net785 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\] _0713_ _0606_
+ VPWR VGND sg13g2_mux2_1
X_4899__52 VPWR VGND net52 sg13g2_tiehi
X_4407_ _2051_ _2048_ _2050_ VPWR VGND sg13g2_xnor2_1
X_2599_ VPWR _0655_ tmds_blue.dc_balancing_reg\[4\] VGND sg13g2_inv_1
X_4338_ _0914_ net606 _1991_ VPWR VGND sg13g2_nor2b_1
X_4269_ _1913_ _1923_ _1924_ _1930_ _1931_ VPWR VGND sg13g2_and4_1
XFILLER_15_506 VPWR VGND sg13g2_fill_1
XFILLER_15_528 VPWR VGND sg13g2_decap_4
XFILLER_42_347 VPWR VGND sg13g2_decap_8
XFILLER_11_734 VPWR VGND sg13g2_decap_4
XFILLER_10_211 VPWR VGND sg13g2_fill_2
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_11_789 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_fill_1
XFILLER_6_259 VPWR VGND sg13g2_decap_8
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_46_1021 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
Xfanout780 net783 net780 VPWR VGND sg13g2_buf_8
XFILLER_18_311 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_fill_1
XFILLER_45_163 VPWR VGND sg13g2_decap_4
XFILLER_42_892 VPWR VGND sg13g2_decap_8
X_5119__213 VPWR VGND net213 sg13g2_tiehi
X_3640_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\] net569 _1309_ VPWR
+ VGND sg13g2_nor2_1
X_3571_ _1213_ _1219_ _1239_ _1240_ VPWR VGND sg13g2_or3_1
XFILLER_6_771 VPWR VGND sg13g2_fill_1
X_5241_ net802 VGND VPWR serialize.n427\[2\] serialize.n411\[0\] clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_5_292 VPWR VGND sg13g2_decap_8
X_5172_ net132 VGND VPWR _0596_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[2\]
+ _0244_ sg13g2_dfrbpq_1
X_4123_ _1294_ _1779_ _1787_ _1788_ VPWR VGND sg13g2_nor3_1
X_4054_ VPWR VGND _1716_ _1718_ _1715_ _1711_ _1719_ _1712_ sg13g2_a221oi_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_2
X_3005_ net779 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\] _0803_ _0268_
+ VPWR VGND sg13g2_mux2_1
XFILLER_24_314 VPWR VGND sg13g2_decap_8
X_5102__283 VPWR VGND net283 sg13g2_tiehi
X_4956_ net328 VGND VPWR _0384_ red_tmds_par\[2\] net641 sg13g2_dfrbpq_1
X_4887_ net75 VGND VPWR _0315_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\]
+ _0036_ sg13g2_dfrbpq_1
XFILLER_20_531 VPWR VGND sg13g2_fill_2
X_3907_ net616 _1570_ _1575_ _1576_ VPWR VGND sg13g2_nor3_1
XFILLER_32_380 VPWR VGND sg13g2_fill_1
X_3838_ net622 _1501_ _1506_ _1507_ VPWR VGND sg13g2_nor3_1
XFILLER_4_708 VPWR VGND sg13g2_decap_4
XFILLER_4_719 VPWR VGND sg13g2_fill_1
X_3769_ _1434_ _1435_ _1436_ _1437_ _1438_ VPWR VGND sg13g2_nor4_1
XFILLER_10_34 VPWR VGND sg13g2_decap_4
XFILLER_10_78 VPWR VGND sg13g2_fill_1
XFILLER_0_936 VPWR VGND sg13g2_decap_8
XFILLER_48_907 VPWR VGND sg13g2_decap_8
XFILLER_19_21 VPWR VGND sg13g2_decap_4
XFILLER_19_108 VPWR VGND sg13g2_fill_2
XFILLER_28_620 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_4
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_24_892 VPWR VGND sg13g2_decap_8
XFILLER_11_575 VPWR VGND sg13g2_decap_4
X_5188__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_2_273 VPWR VGND sg13g2_fill_1
XFILLER_19_631 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_46_450 VPWR VGND sg13g2_decap_8
XFILLER_19_653 VPWR VGND sg13g2_fill_2
XFILLER_46_494 VPWR VGND sg13g2_decap_4
XFILLER_33_111 VPWR VGND sg13g2_decap_8
XFILLER_34_656 VPWR VGND sg13g2_decap_8
X_4810_ net688 net740 _0240_ VPWR VGND sg13g2_nor2_1
XFILLER_21_306 VPWR VGND sg13g2_decap_4
XFILLER_33_155 VPWR VGND sg13g2_decap_4
X_4741_ net656 net708 _0171_ VPWR VGND sg13g2_nor2_1
X_4672_ net685 net737 _0102_ VPWR VGND sg13g2_nor2_1
X_3623_ VGND VPWR _1290_ _1291_ _1292_ _1282_ sg13g2_a21oi_1
X_3554_ _1213_ _1066_ _1223_ VPWR VGND _1218_ sg13g2_nand3b_1
X_3485_ _1098_ _1143_ _1097_ _1154_ VPWR VGND sg13g2_nand3_1
X_5224_ net804 VGND VPWR net420 serialize.n420\[4\] clknet_3_2__leaf_clk_regs sg13g2_dfrbpq_1
X_5155_ net289 VGND VPWR _0579_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\]
+ _0227_ sg13g2_dfrbpq_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_4106_ _1703_ _1754_ _1771_ VPWR VGND sg13g2_nor2_1
X_5086_ net361 VGND VPWR _0510_ tmds_red.dc_balancing_reg\[1\] net644 sg13g2_dfrbpq_2
X_4037_ _0990_ VPWR _1702_ VGND _0989_ _1059_ sg13g2_o21ai_1
X_5026__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_24_100 VPWR VGND sg13g2_decap_4
XFILLER_12_328 VPWR VGND sg13g2_decap_4
X_4939_ net345 VGND VPWR _0367_ videogen.test_lut_thingy.gol_counter_reg\[1\] net639
+ sg13g2_dfrbpq_2
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_44 VPWR VGND sg13g2_decap_4
X_4911__400 VPWR VGND net400 sg13g2_tiehi
XFILLER_0_733 VPWR VGND sg13g2_decap_8
XFILLER_48_715 VPWR VGND sg13g2_fill_1
X_4983__280 VPWR VGND net280 sg13g2_tiehi
XFILLER_29_951 VPWR VGND sg13g2_decap_8
XFILLER_44_943 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_fill_1
XFILLER_43_442 VPWR VGND sg13g2_fill_1
XFILLER_15_133 VPWR VGND sg13g2_fill_1
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_8_877 VPWR VGND sg13g2_decap_8
XFILLER_7_68 VPWR VGND sg13g2_decap_8
X_3270_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\] _0968_ _0971_ VPWR
+ VGND sg13g2_and2_1
XFILLER_46_280 VPWR VGND sg13g2_fill_2
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_21_103 VPWR VGND sg13g2_fill_1
XFILLER_21_114 VPWR VGND sg13g2_decap_8
X_4724_ net650 net703 _0154_ VPWR VGND sg13g2_nor2_1
X_2985_ net773 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\] _0799_ _0292_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_681 VPWR VGND sg13g2_decap_8
X_4655_ net670 net721 _0085_ VPWR VGND sg13g2_nor2_1
X_4586_ net657 net709 _0016_ VPWR VGND sg13g2_nor2_1
X_3606_ _1273_ _1274_ _1275_ VPWR VGND sg13g2_nor2_1
XFILLER_1_508 VPWR VGND sg13g2_decap_8
X_3537_ _1203_ _1204_ _1198_ _1206_ VPWR VGND sg13g2_nand3_1
XFILLER_27_1019 VPWR VGND sg13g2_decap_8
X_3468_ _1113_ _1130_ _1112_ _1137_ VPWR VGND _1131_ sg13g2_nand4_1
X_5207_ net403 VGND VPWR _0631_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\]
+ _0261_ sg13g2_dfrbpq_1
X_3399_ VPWR VGND _0993_ _0992_ _0991_ videogen.fancy_shader.video_y\[3\] _1068_ videogen.fancy_shader.n646\[3\]
+ sg13g2_a221oi_1
XFILLER_29_203 VPWR VGND sg13g2_decap_4
X_5180__347 VPWR VGND net347 sg13g2_tiehi
XFILLER_29_225 VPWR VGND sg13g2_decap_4
X_5138_ net104 VGND VPWR _0562_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\]
+ _0210_ sg13g2_dfrbpq_1
XFILLER_29_269 VPWR VGND sg13g2_decap_8
X_5069_ net47 VGND VPWR _0493_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\]
+ _0150_ sg13g2_dfrbpq_1
XFILLER_26_965 VPWR VGND sg13g2_decap_8
XFILLER_13_626 VPWR VGND sg13g2_fill_1
XFILLER_16_77 VPWR VGND sg13g2_decap_4
XFILLER_25_475 VPWR VGND sg13g2_fill_2
XFILLER_40_434 VPWR VGND sg13g2_decap_4
XFILLER_9_608 VPWR VGND sg13g2_fill_2
XFILLER_12_136 VPWR VGND sg13g2_decap_4
XFILLER_13_637 VPWR VGND sg13g2_fill_2
XFILLER_41_979 VPWR VGND sg13g2_decap_8
XFILLER_40_489 VPWR VGND sg13g2_decap_8
XFILLER_20_191 VPWR VGND sg13g2_fill_2
XFILLER_5_847 VPWR VGND sg13g2_decap_4
XFILLER_4_324 VPWR VGND sg13g2_decap_8
XFILLER_4_302 VPWR VGND sg13g2_decap_8
XFILLER_48_545 VPWR VGND sg13g2_decap_8
XFILLER_17_954 VPWR VGND sg13g2_decap_8
XFILLER_44_773 VPWR VGND sg13g2_fill_1
XFILLER_43_294 VPWR VGND sg13g2_fill_2
XFILLER_31_434 VPWR VGND sg13g2_decap_8
XFILLER_32_957 VPWR VGND sg13g2_decap_8
XFILLER_31_478 VPWR VGND sg13g2_decap_4
X_2770_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\] _0746_ _0537_
+ VPWR VGND sg13g2_mux2_1
X_4440_ _0618_ _2076_ net572 _2070_ net607 VPWR VGND sg13g2_a22oi_1
X_4371_ _2017_ net548 _1996_ VPWR VGND sg13g2_nand2_1
Xfanout609 videogen.fancy_shader.n646\[8\] net609 VPWR VGND sg13g2_buf_8
X_3322_ _1006_ _1002_ _1012_ VPWR VGND sg13g2_xor2_1
X_3253_ VGND VPWR net628 _0957_ _0960_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\]
+ sg13g2_a21oi_1
X_3184_ _0906_ net547 _0913_ VPWR VGND sg13g2_nor2b_2
XFILLER_23_902 VPWR VGND sg13g2_decap_8
XFILLER_23_979 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
X_2968_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\] _0794_ _0314_
+ VPWR VGND sg13g2_mux2_1
X_4707_ net651 net701 _0137_ VPWR VGND sg13g2_nor2_1
X_4638_ net663 net716 _0068_ VPWR VGND sg13g2_nor2_1
X_2899_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\] net777 _0777_ _0430_
+ VPWR VGND sg13g2_mux2_1
X_4569_ _2197_ _2194_ _2196_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_817 VPWR VGND sg13g2_decap_8
XFILLER_49_309 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_45_537 VPWR VGND sg13g2_decap_8
XFILLER_45_526 VPWR VGND sg13g2_fill_2
XFILLER_27_32 VPWR VGND sg13g2_decap_4
XFILLER_27_76 VPWR VGND sg13g2_fill_1
XFILLER_14_924 VPWR VGND sg13g2_decap_8
XFILLER_40_220 VPWR VGND sg13g2_fill_1
XFILLER_9_416 VPWR VGND sg13g2_fill_1
XFILLER_13_467 VPWR VGND sg13g2_decap_8
XFILLER_5_666 VPWR VGND sg13g2_fill_2
XFILLER_4_187 VPWR VGND sg13g2_fill_1
XFILLER_4_69 VPWR VGND sg13g2_decap_8
XFILLER_1_872 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_8
XFILLER_48_353 VPWR VGND sg13g2_decap_8
XFILLER_17_751 VPWR VGND sg13g2_decap_8
X_3940_ net625 VPWR _1608_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\]
+ net590 sg13g2_o21ai_1
X_3871_ VGND VPWR _1533_ _1539_ _1540_ net611 sg13g2_a21oi_1
X_2822_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\] net780 _0756_ _0486_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_927 VPWR VGND sg13g2_decap_8
XFILLER_32_787 VPWR VGND sg13g2_fill_2
X_2753_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\] net765 _0740_ _0548_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
X_2684_ net792 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\] _0721_ _0598_
+ VPWR VGND sg13g2_mux2_1
X_4423_ _2065_ tmds_blue.n193 net603 VPWR VGND sg13g2_nand2b_1
X_4354_ VPWR _2000_ _1999_ VGND sg13g2_inv_1
X_3305_ net750 _0984_ _0996_ _0348_ VPWR VGND sg13g2_nor3_1
X_4285_ _1936_ _1946_ _1947_ VPWR VGND sg13g2_nor2_1
X_3236_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0946_ _0948_ VPWR VGND
+ sg13g2_and2_1
X_5064__262 VPWR VGND net262 sg13g2_tiehi
X_3167_ _0895_ VPWR _0896_ VGND _0883_ _0893_ sg13g2_o21ai_1
XFILLER_27_526 VPWR VGND sg13g2_decap_8
X_3098_ net429 green_tmds_par\[6\] net695 serialize.n428\[6\] VPWR VGND sg13g2_mux2_1
XFILLER_14_209 VPWR VGND sg13g2_fill_1
XFILLER_23_743 VPWR VGND sg13g2_fill_2
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_23_798 VPWR VGND sg13g2_fill_1
XFILLER_2_614 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_4
XFILLER_49_128 VPWR VGND sg13g2_decap_8
XFILLER_45_312 VPWR VGND sg13g2_fill_2
XFILLER_46_846 VPWR VGND sg13g2_decap_8
XFILLER_41_562 VPWR VGND sg13g2_fill_2
XFILLER_14_798 VPWR VGND sg13g2_decap_4
XFILLER_6_942 VPWR VGND sg13g2_decap_8
XFILLER_10_993 VPWR VGND sg13g2_decap_8
X_4070_ _1735_ _1717_ _1724_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_1000 VPWR VGND sg13g2_decap_8
X_3021_ _0651_ _0680_ _0817_ VPWR VGND sg13g2_and2_1
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_48_183 VPWR VGND sg13g2_fill_1
XFILLER_48_172 VPWR VGND sg13g2_decap_8
X_4972_ net301 VGND VPWR _0400_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\]
+ _0057_ sg13g2_dfrbpq_1
X_3923_ net749 net1 _1592_ VPWR VGND sg13g2_nor2_1
X_4959__325 VPWR VGND net325 sg13g2_tiehi
X_3854_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\] net588 _1523_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_713 VPWR VGND sg13g2_decap_4
XFILLER_32_584 VPWR VGND sg13g2_fill_1
X_2805_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\] net753 _0753_ _0500_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_735 VPWR VGND sg13g2_decap_4
X_3785_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\] net590 _1454_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
X_2736_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\] _0736_ _0561_
+ VPWR VGND sg13g2_mux2_1
X_2667_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\] _0713_ _0607_
+ VPWR VGND sg13g2_mux2_1
X_4902__46 VPWR VGND net46 sg13g2_tiehi
X_4406_ _2050_ _0664_ _2049_ VPWR VGND sg13g2_xnor2_1
X_2598_ tmds_green.dc_balancing_reg\[4\] _0654_ VPWR VGND sg13g2_inv_4
X_4337_ net749 _1990_ _0387_ VPWR VGND sg13g2_nor2_1
X_4268_ _1930_ _1928_ _1929_ VPWR VGND sg13g2_nand2_1
X_3219_ _0923_ _0934_ _0308_ VPWR VGND sg13g2_nor2_1
X_4199_ _1856_ _1859_ _1855_ _1861_ VPWR VGND sg13g2_nand3_1
XFILLER_27_323 VPWR VGND sg13g2_fill_1
XFILLER_15_518 VPWR VGND sg13g2_decap_4
XFILLER_27_367 VPWR VGND sg13g2_decap_8
XFILLER_28_879 VPWR VGND sg13g2_fill_1
XFILLER_27_389 VPWR VGND sg13g2_fill_1
XFILLER_23_551 VPWR VGND sg13g2_fill_2
XFILLER_10_234 VPWR VGND sg13g2_fill_1
XFILLER_6_238 VPWR VGND sg13g2_decap_8
X_5036__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_40_87 VPWR VGND sg13g2_fill_1
XFILLER_46_1000 VPWR VGND sg13g2_decap_8
XFILLER_3_934 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
Xfanout770 net771 net770 VPWR VGND sg13g2_buf_8
Xfanout781 net783 net781 VPWR VGND sg13g2_buf_8
Xfanout792 net793 net792 VPWR VGND sg13g2_buf_8
XFILLER_45_142 VPWR VGND sg13g2_decap_8
XFILLER_18_356 VPWR VGND sg13g2_fill_1
XFILLER_34_816 VPWR VGND sg13g2_fill_2
XFILLER_45_175 VPWR VGND sg13g2_fill_1
XFILLER_33_315 VPWR VGND sg13g2_decap_8
XFILLER_42_871 VPWR VGND sg13g2_fill_1
XFILLER_42_860 VPWR VGND sg13g2_decap_8
XFILLER_14_584 VPWR VGND sg13g2_decap_8
XFILLER_14_595 VPWR VGND sg13g2_fill_1
X_3570_ VPWR VGND _1230_ _1220_ _1227_ _1061_ _1239_ _1062_ sg13g2_a221oi_1
X_5240_ net805 VGND VPWR serialize.n427\[1\] serialize.n452 clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_5_260 VPWR VGND sg13g2_fill_2
X_5171_ net159 VGND VPWR _0595_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[1\]
+ _0243_ sg13g2_dfrbpq_1
X_4122_ _1767_ _1772_ _1787_ VPWR VGND sg13g2_and2_1
X_4053_ _1718_ _1147_ _1709_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_481 VPWR VGND sg13g2_decap_4
X_3004_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\] _0803_ _0269_
+ VPWR VGND sg13g2_mux2_1
X_5096__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_24_359 VPWR VGND sg13g2_decap_8
X_4955_ net329 VGND VPWR _0383_ tmds_red.n132 net642 sg13g2_dfrbpq_2
X_3906_ net626 _1571_ _1572_ _1574_ _1575_ VPWR VGND sg13g2_nor4_1
XFILLER_33_893 VPWR VGND sg13g2_decap_4
X_4886_ net77 VGND VPWR _0314_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\]
+ _0035_ sg13g2_dfrbpq_1
X_3837_ _1502_ _1503_ _1504_ _1505_ _1506_ VPWR VGND sg13g2_nor4_1
XFILLER_20_565 VPWR VGND sg13g2_decap_4
X_3768_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\] net574 _1437_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_598 VPWR VGND sg13g2_decap_8
X_2719_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\] _0731_ _0573_
+ VPWR VGND sg13g2_mux2_1
XFILLER_3_219 VPWR VGND sg13g2_fill_2
X_3699_ VGND VPWR _0634_ net593 _1368_ _1367_ sg13g2_a21oi_1
XFILLER_0_915 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_28_665 VPWR VGND sg13g2_decap_4
XFILLER_28_676 VPWR VGND sg13g2_decap_4
XFILLER_43_635 VPWR VGND sg13g2_decap_4
XFILLER_43_613 VPWR VGND sg13g2_fill_1
XFILLER_15_315 VPWR VGND sg13g2_fill_1
XFILLER_27_164 VPWR VGND sg13g2_fill_2
XFILLER_28_698 VPWR VGND sg13g2_fill_2
XFILLER_35_54 VPWR VGND sg13g2_fill_2
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_23_381 VPWR VGND sg13g2_fill_2
XFILLER_7_514 VPWR VGND sg13g2_fill_2
XFILLER_7_503 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_4
XFILLER_11_554 VPWR VGND sg13g2_decap_8
XFILLER_13_1010 VPWR VGND sg13g2_decap_8
XFILLER_7_558 VPWR VGND sg13g2_decap_8
XFILLER_7_536 VPWR VGND sg13g2_decap_4
XFILLER_2_252 VPWR VGND sg13g2_decap_8
XFILLER_2_285 VPWR VGND sg13g2_fill_2
X_4949__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_38_407 VPWR VGND sg13g2_fill_1
XFILLER_38_418 VPWR VGND sg13g2_decap_4
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_19_665 VPWR VGND sg13g2_decap_4
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_21_318 VPWR VGND sg13g2_fill_2
X_4740_ net656 net711 _0170_ VPWR VGND sg13g2_nor2_1
XFILLER_33_189 VPWR VGND sg13g2_decap_4
X_4956__328 VPWR VGND net328 sg13g2_tiehi
X_4671_ net653 net705 _0101_ VPWR VGND sg13g2_nor2_1
XFILLER_30_852 VPWR VGND sg13g2_fill_2
XFILLER_30_874 VPWR VGND sg13g2_decap_4
X_3622_ VGND VPWR _1276_ _1279_ _1291_ _1235_ sg13g2_a21oi_1
X_3553_ VGND VPWR _1222_ _1221_ _1220_ sg13g2_or2_1
XFILLER_44_0 VPWR VGND sg13g2_decap_4
X_3484_ _1143_ _1098_ _1096_ _1153_ VPWR VGND sg13g2_a21o_1
X_5223_ net804 VGND VPWR serialize.n431\[5\] serialize.n420\[3\] clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5154_ net297 VGND VPWR _0578_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\]
+ _0226_ sg13g2_dfrbpq_1
X_4105_ _1770_ _1769_ _1768_ VPWR VGND sg13g2_nand2b_1
X_5085_ net363 VGND VPWR _0509_ tmds_red.dc_balancing_reg\[0\] net644 sg13g2_dfrbpq_1
X_4036_ _1298_ net798 _1701_ _0375_ VPWR VGND sg13g2_a21o_1
XFILLER_21_830 VPWR VGND sg13g2_decap_4
X_4938_ net346 VGND VPWR _0366_ videogen.test_lut_thingy.gol_counter_reg\[0\] net639
+ sg13g2_dfrbpq_2
XFILLER_21_874 VPWR VGND sg13g2_fill_1
X_4869_ net101 VGND VPWR _0297_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\]
+ _0028_ sg13g2_dfrbpq_1
XFILLER_21_89 VPWR VGND sg13g2_decap_8
XFILLER_0_712 VPWR VGND sg13g2_decap_8
XFILLER_43_1025 VPWR VGND sg13g2_decap_4
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_29_930 VPWR VGND sg13g2_decap_8
XFILLER_44_922 VPWR VGND sg13g2_decap_8
XFILLER_16_646 VPWR VGND sg13g2_decap_8
XFILLER_16_657 VPWR VGND sg13g2_fill_2
XFILLER_44_999 VPWR VGND sg13g2_decap_8
XFILLER_43_487 VPWR VGND sg13g2_fill_1
XFILLER_43_465 VPWR VGND sg13g2_decap_8
XFILLER_43_454 VPWR VGND sg13g2_fill_2
XFILLER_16_679 VPWR VGND sg13g2_fill_2
XFILLER_31_616 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_4
XFILLER_30_148 VPWR VGND sg13g2_fill_1
XFILLER_7_300 VPWR VGND sg13g2_decap_8
XFILLER_3_550 VPWR VGND sg13g2_fill_1
XFILLER_3_583 VPWR VGND sg13g2_decap_4
XFILLER_16_4 VPWR VGND sg13g2_decap_4
XFILLER_38_259 VPWR VGND sg13g2_fill_1
X_4962__321 VPWR VGND net321 sg13g2_tiehi
XFILLER_35_955 VPWR VGND sg13g2_decap_8
XFILLER_34_476 VPWR VGND sg13g2_decap_4
X_2984_ net762 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\] _0799_ _0293_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_690 VPWR VGND sg13g2_fill_1
X_4723_ net655 net707 _0153_ VPWR VGND sg13g2_nor2_1
X_4654_ net670 net721 _0084_ VPWR VGND sg13g2_nor2_1
X_3605_ _1196_ _1271_ _1274_ VPWR VGND sg13g2_and2_1
X_4585_ net652 net704 _0015_ VPWR VGND sg13g2_nor2_1
X_3536_ _1205_ _1203_ _1204_ VPWR VGND sg13g2_nand2_1
X_3467_ _1136_ _1132_ _1133_ _1111_ _1110_ VPWR VGND sg13g2_a22oi_1
X_5206_ net250 VGND VPWR _0630_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\]
+ _0260_ sg13g2_dfrbpq_1
X_3398_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.n646\[3\] _1067_
+ VPWR VGND sg13g2_nor2_1
X_5137_ net112 VGND VPWR _0561_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\]
+ _0209_ sg13g2_dfrbpq_1
X_5068_ net51 VGND VPWR _0001_ videogen.test_lut_thingy.pixel_feeder_inst.state\[3\]
+ net635 sg13g2_dfrbpq_1
X_4019_ _1686_ VPWR _1687_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\]
+ net588 sg13g2_o21ai_1
XFILLER_37_292 VPWR VGND sg13g2_decap_4
XFILLER_25_410 VPWR VGND sg13g2_decap_8
XFILLER_25_443 VPWR VGND sg13g2_decap_8
XFILLER_26_944 VPWR VGND sg13g2_decap_8
XFILLER_16_45 VPWR VGND sg13g2_decap_4
XFILLER_12_115 VPWR VGND sg13g2_fill_2
X_4939__345 VPWR VGND net345 sg13g2_tiehi
XFILLER_21_693 VPWR VGND sg13g2_fill_2
XFILLER_4_369 VPWR VGND sg13g2_decap_8
XFILLER_0_564 VPWR VGND sg13g2_decap_8
XFILLER_48_524 VPWR VGND sg13g2_decap_8
X_4946__338 VPWR VGND net338 sg13g2_tiehi
XFILLER_44_741 VPWR VGND sg13g2_fill_1
XFILLER_17_933 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_16_487 VPWR VGND sg13g2_decap_4
XFILLER_32_936 VPWR VGND sg13g2_decap_8
XFILLER_11_170 VPWR VGND sg13g2_decap_4
X_4370_ _2016_ _2014_ _2015_ _2008_ _0913_ VPWR VGND sg13g2_a22oi_1
X_3321_ _1005_ _1010_ _1011_ VPWR VGND sg13g2_nor2_2
X_3252_ net578 _0956_ _0959_ VPWR VGND sg13g2_nor2_1
XFILLER_39_524 VPWR VGND sg13g2_decap_8
X_3183_ VPWR _0912_ _0911_ VGND sg13g2_inv_1
X_5197__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_26_218 VPWR VGND sg13g2_fill_1
XFILLER_22_402 VPWR VGND sg13g2_decap_4
XFILLER_23_958 VPWR VGND sg13g2_decap_8
X_2967_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\] _0794_ _0315_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_991 VPWR VGND sg13g2_decap_8
X_4706_ net652 net704 _0136_ VPWR VGND sg13g2_nor2_1
X_5134__136 VPWR VGND net136 sg13g2_tiehi
X_2898_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\] net764 _0777_ _0431_
+ VPWR VGND sg13g2_mux2_1
X_4637_ net664 net715 _0067_ VPWR VGND sg13g2_nor2_1
X_4568_ _2196_ _0655_ _2195_ VPWR VGND sg13g2_xnor2_1
X_4499_ _0856_ _2122_ _2131_ _2132_ VPWR VGND sg13g2_nor3_1
X_3519_ _1184_ _1186_ _1077_ _1188_ VPWR VGND sg13g2_nand3_1
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
XFILLER_18_719 VPWR VGND sg13g2_fill_2
XFILLER_38_590 VPWR VGND sg13g2_fill_1
XFILLER_14_903 VPWR VGND sg13g2_decap_8
XFILLER_13_402 VPWR VGND sg13g2_decap_4
XFILLER_13_424 VPWR VGND sg13g2_fill_2
XFILLER_26_785 VPWR VGND sg13g2_decap_4
XFILLER_43_54 VPWR VGND sg13g2_fill_1
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_4_15 VPWR VGND sg13g2_fill_2
XFILLER_4_59 VPWR VGND sg13g2_decap_4
XFILLER_1_851 VPWR VGND sg13g2_decap_8
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_0_383 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_fill_1
XFILLER_32_733 VPWR VGND sg13g2_decap_8
X_3870_ net624 _1538_ _1539_ VPWR VGND sg13g2_nor2_1
XFILLER_20_906 VPWR VGND sg13g2_decap_8
X_2821_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\] net768 _0756_ _0487_
+ VPWR VGND sg13g2_mux2_1
X_2752_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\] net756 _0740_ _0549_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_298 VPWR VGND sg13g2_fill_2
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_4422_ VGND VPWR net605 _2063_ _0610_ _2064_ sg13g2_a21oi_1
X_2683_ net782 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[1\] _0721_ _0599_
+ VPWR VGND sg13g2_mux2_1
X_4353_ _1999_ tmds_red.dc_balancing_reg\[2\] _0905_ VPWR VGND sg13g2_xnor2_1
X_3304_ _0942_ _0995_ _0996_ VPWR VGND sg13g2_nor2b_2
X_4284_ _1931_ _1940_ _1946_ VPWR VGND sg13g2_nor2_1
X_3235_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0946_ _0947_ VPWR VGND
+ sg13g2_nor2_1
X_3166_ _0895_ _0883_ _0894_ VPWR VGND sg13g2_nand2_1
X_3097_ _0850_ VPWR serialize.n428\[5\] VGND _0670_ net698 sg13g2_o21ai_1
XFILLER_27_549 VPWR VGND sg13g2_fill_1
XFILLER_42_508 VPWR VGND sg13g2_fill_2
X_5105__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_35_593 VPWR VGND sg13g2_decap_4
X_3999_ VGND VPWR _1667_ _1666_ _1655_ sg13g2_or2_1
XFILLER_11_917 VPWR VGND sg13g2_decap_8
XFILLER_22_254 VPWR VGND sg13g2_decap_8
XFILLER_6_409 VPWR VGND sg13g2_fill_1
XFILLER_13_68 VPWR VGND sg13g2_decap_8
XFILLER_2_604 VPWR VGND sg13g2_fill_1
XFILLER_2_637 VPWR VGND sg13g2_fill_2
XFILLER_14_722 VPWR VGND sg13g2_fill_1
XFILLER_26_560 VPWR VGND sg13g2_decap_8
XFILLER_13_232 VPWR VGND sg13g2_fill_1
XFILLER_13_276 VPWR VGND sg13g2_decap_8
XFILLER_9_236 VPWR VGND sg13g2_fill_2
XFILLER_13_298 VPWR VGND sg13g2_fill_1
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_10_972 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_497 VPWR VGND sg13g2_decap_8
XFILLER_49_674 VPWR VGND sg13g2_fill_2
X_3020_ videogen.fancy_shader.video_x\[6\] _0815_ _0816_ VPWR VGND sg13g2_and2_1
XFILLER_48_195 VPWR VGND sg13g2_decap_8
XFILLER_37_858 VPWR VGND sg13g2_decap_4
XFILLER_17_571 VPWR VGND sg13g2_fill_2
X_4971_ net303 VGND VPWR _0399_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[2\]
+ _0056_ sg13g2_dfrbpq_1
X_3922_ _1591_ _1542_ _1590_ videogen.test_lut_thingy.gol_counter_reg\[3\] _0661_
+ VPWR VGND sg13g2_a22oi_1
X_3853_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\] net557 _1522_ VPWR
+ VGND sg13g2_nor2_1
X_2804_ _0700_ _0737_ _0753_ VPWR VGND sg13g2_nor2_2
X_3784_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\] net568 _1453_ VPWR
+ VGND sg13g2_nor2_1
X_2735_ _0736_ _0711_ _0732_ VPWR VGND sg13g2_nand2_2
X_2666_ net763 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\] _0713_ _0608_
+ VPWR VGND sg13g2_mux2_1
X_4405_ VGND VPWR tmds_red.dc_balancing_reg\[3\] _2023_ _2049_ _0902_ sg13g2_a21oi_1
X_2597_ VPWR _0653_ tmds_green.dc_balancing_reg\[3\] VGND sg13g2_inv_1
X_4336_ net547 net607 _1990_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
X_4267_ _1929_ _1800_ _1927_ VPWR VGND sg13g2_nand2_1
X_4849__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_39_140 VPWR VGND sg13g2_decap_8
X_3218_ _0932_ videogen.fancy_shader.video_x\[9\] _0934_ VPWR VGND sg13g2_xor2_1
X_4198_ VPWR _1860_ _1859_ VGND sg13g2_inv_1
XFILLER_27_302 VPWR VGND sg13g2_fill_1
XFILLER_28_803 VPWR VGND sg13g2_decap_8
XFILLER_28_814 VPWR VGND sg13g2_fill_2
X_3149_ _0878_ _0876_ _0877_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_213 VPWR VGND sg13g2_fill_1
XFILLER_24_78 VPWR VGND sg13g2_decap_4
XFILLER_3_913 VPWR VGND sg13g2_decap_8
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
Xfanout760 net761 net760 VPWR VGND sg13g2_buf_8
Xfanout771 net772 net771 VPWR VGND sg13g2_buf_8
Xfanout793 net794 net793 VPWR VGND sg13g2_buf_8
Xfanout782 net783 net782 VPWR VGND sg13g2_buf_8
XFILLER_18_368 VPWR VGND sg13g2_fill_2
XFILLER_19_869 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_4
XFILLER_33_327 VPWR VGND sg13g2_fill_2
X_5170_ net167 VGND VPWR _0594_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\]
+ _0242_ sg13g2_dfrbpq_1
X_4121_ _1770_ VPWR _1786_ VGND _1703_ _1777_ sg13g2_o21ai_1
X_4052_ _1717_ _1715_ _1716_ VPWR VGND sg13g2_nand2_2
X_3003_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\] _0803_ _0270_
+ VPWR VGND sg13g2_mux2_1
X_5058__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_37_699 VPWR VGND sg13g2_decap_8
XFILLER_25_828 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_fill_2
X_4954_ net330 VGND VPWR _0382_ tmds_red.n126 net642 sg13g2_dfrbpq_2
X_3905_ _1573_ VPWR _1574_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[3\]
+ net569 sg13g2_o21ai_1
X_4885_ net79 VGND VPWR _0313_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[0\]
+ _0034_ sg13g2_dfrbpq_1
X_3836_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\] net568 _1505_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_544 VPWR VGND sg13g2_decap_8
X_4972__301 VPWR VGND net301 sg13g2_tiehi
X_3767_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\] net551 _1436_ VPWR
+ VGND sg13g2_nor2_1
X_2718_ _0731_ _0716_ VPWR VGND _0719_ sg13g2_nand2b_2
X_3698_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\] net553 _1367_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_10_69 VPWR VGND sg13g2_decap_8
XFILLER_10_58 VPWR VGND sg13g2_decap_8
X_2649_ _0702_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\] net628 VPWR VGND
+ sg13g2_nand2_2
X_4319_ _1978_ _1974_ _1977_ _1698_ _1593_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_132 VPWR VGND sg13g2_decap_4
XFILLER_27_187 VPWR VGND sg13g2_decap_8
XFILLER_2_220 VPWR VGND sg13g2_fill_1
XFILLER_2_231 VPWR VGND sg13g2_decap_4
XFILLER_3_787 VPWR VGND sg13g2_decap_8
X_5142__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_47_920 VPWR VGND sg13g2_decap_8
Xfanout590 net592 net590 VPWR VGND sg13g2_buf_8
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
XFILLER_19_655 VPWR VGND sg13g2_fill_1
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_34_647 VPWR VGND sg13g2_decap_4
XFILLER_15_861 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_fill_2
X_4670_ net653 net706 _0100_ VPWR VGND sg13g2_nor2_1
X_3621_ _1278_ _1065_ _1275_ _1290_ VPWR VGND sg13g2_a21o_1
X_3552_ _1221_ _1064_ _1213_ VPWR VGND sg13g2_nand2_1
X_3483_ _1098_ _1143_ _1096_ _1152_ VPWR VGND sg13g2_nand3_1
X_5222_ net804 VGND VPWR serialize.n431\[4\] serialize.n420\[2\] clknet_3_3__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5153_ net304 VGND VPWR _0577_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\]
+ _0225_ sg13g2_dfrbpq_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_4104_ _1762_ _1765_ _1757_ _1769_ VPWR VGND sg13g2_nand3_1
X_5084_ net365 VGND VPWR _0508_ green_tmds_par\[9\] net646 sg13g2_dfrbpq_1
XFILLER_49_290 VPWR VGND sg13g2_decap_8
X_4035_ VGND VPWR _1398_ _1700_ _1701_ _1594_ sg13g2_a21oi_1
XFILLER_38_986 VPWR VGND sg13g2_decap_8
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_fill_1
X_4937_ net348 VGND VPWR _0365_ videogen.fancy_shader.video_y\[9\] net632 sg13g2_dfrbpq_2
X_5137__112 VPWR VGND net112 sg13g2_tiehi
X_4868_ net103 VGND VPWR _0296_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[1\]
+ _0027_ sg13g2_dfrbpq_1
X_3819_ _1486_ VPWR _1488_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\]
+ net556 sg13g2_o21ai_1
X_4799_ net691 net742 _0229_ VPWR VGND sg13g2_nor2_1
XFILLER_43_1004 VPWR VGND sg13g2_decap_8
XFILLER_0_768 VPWR VGND sg13g2_decap_8
XFILLER_47_249 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_4
X_5005__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_43_422 VPWR VGND sg13g2_fill_2
XFILLER_28_496 VPWR VGND sg13g2_decap_8
XFILLER_44_978 VPWR VGND sg13g2_decap_8
X_5079__379 VPWR VGND net379 sg13g2_tiehi
XFILLER_8_813 VPWR VGND sg13g2_fill_2
X_5155__289 VPWR VGND net289 sg13g2_tiehi
XFILLER_7_356 VPWR VGND sg13g2_fill_2
XFILLER_7_345 VPWR VGND sg13g2_decap_8
XFILLER_3_562 VPWR VGND sg13g2_decap_8
XFILLER_11_90 VPWR VGND sg13g2_decap_8
XFILLER_3_595 VPWR VGND sg13g2_fill_1
XFILLER_39_706 VPWR VGND sg13g2_fill_2
X_2983_ net753 videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\] _0799_ _0294_
+ VPWR VGND sg13g2_mux2_1
X_4722_ net656 net707 _0152_ VPWR VGND sg13g2_nor2_1
X_4653_ net671 net721 _0083_ VPWR VGND sg13g2_nor2_1
X_3604_ _1195_ _1272_ _1273_ VPWR VGND sg13g2_and2_1
X_4584_ net652 net704 _0014_ VPWR VGND sg13g2_nor2_1
X_4852__135 VPWR VGND net135 sg13g2_tiehi
X_3535_ _1170_ VPWR _1204_ VGND _1177_ _1202_ sg13g2_o21ai_1
X_3466_ _1111_ _1132_ _1110_ _1135_ VPWR VGND _1133_ sg13g2_nand4_1
X_5205_ net285 VGND VPWR _0629_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\]
+ _0259_ sg13g2_dfrbpq_1
X_3397_ _1066_ _1065_ VPWR VGND sg13g2_inv_2
X_5136_ net120 VGND VPWR _0560_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\]
+ _0208_ sg13g2_dfrbpq_1
XFILLER_45_709 VPWR VGND sg13g2_fill_2
X_5067_ net402 VGND VPWR _0000_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\]
+ net635 sg13g2_dfrbpq_2
X_4018_ _1686_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_26_923 VPWR VGND sg13g2_decap_8
XFILLER_41_915 VPWR VGND sg13g2_fill_2
XFILLER_13_617 VPWR VGND sg13g2_decap_8
XFILLER_40_414 VPWR VGND sg13g2_fill_2
XFILLER_13_639 VPWR VGND sg13g2_fill_1
XFILLER_40_458 VPWR VGND sg13g2_decap_8
XFILLER_21_672 VPWR VGND sg13g2_decap_8
XFILLER_32_45 VPWR VGND sg13g2_decap_4
XFILLER_20_193 VPWR VGND sg13g2_fill_1
XFILLER_10_1014 VPWR VGND sg13g2_decap_8
XFILLER_0_543 VPWR VGND sg13g2_decap_8
XFILLER_17_912 VPWR VGND sg13g2_decap_8
XFILLER_29_783 VPWR VGND sg13g2_decap_4
XFILLER_35_219 VPWR VGND sg13g2_decap_4
XFILLER_16_411 VPWR VGND sg13g2_decap_8
XFILLER_17_989 VPWR VGND sg13g2_decap_8
XFILLER_31_414 VPWR VGND sg13g2_decap_8
XFILLER_8_610 VPWR VGND sg13g2_fill_1
XFILLER_40_992 VPWR VGND sg13g2_decap_8
XFILLER_8_654 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_4
XFILLER_7_142 VPWR VGND sg13g2_fill_1
X_3320_ _1010_ videogen.fancy_shader.n646\[0\] videogen.fancy_shader.video_x\[0\]
+ VPWR VGND sg13g2_xnor2_1
X_3251_ VGND VPWR _0647_ _0956_ _0324_ _0958_ sg13g2_a21oi_1
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
X_3182_ _0911_ _0906_ _0910_ VPWR VGND sg13g2_nand2_1
XFILLER_19_282 VPWR VGND sg13g2_decap_4
XFILLER_34_230 VPWR VGND sg13g2_fill_2
XFILLER_22_414 VPWR VGND sg13g2_fill_1
XFILLER_23_937 VPWR VGND sg13g2_decap_8
X_2966_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[3\] _0794_ _0316_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_970 VPWR VGND sg13g2_decap_8
X_4705_ net649 net701 _0135_ VPWR VGND sg13g2_nor2_1
XFILLER_30_491 VPWR VGND sg13g2_decap_8
X_2897_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\] net755 _0777_ _0432_
+ VPWR VGND sg13g2_mux2_1
X_4636_ net664 net716 _0066_ VPWR VGND sg13g2_nor2_1
X_4567_ _2172_ VPWR _2195_ VGND _0657_ _2140_ sg13g2_o21ai_1
X_4498_ VGND VPWR _2125_ _2130_ _2131_ _0863_ sg13g2_a21oi_1
X_3518_ _1186_ _1184_ _1077_ _1187_ VPWR VGND sg13g2_a21o_1
X_3449_ _1118_ videogen.fancy_shader.n646\[7\] net629 VPWR VGND sg13g2_xnor2_1
X_5119_ net213 VGND VPWR _0543_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\]
+ _0191_ sg13g2_dfrbpq_1
XFILLER_45_528 VPWR VGND sg13g2_fill_1
XFILLER_25_230 VPWR VGND sg13g2_decap_8
XFILLER_25_241 VPWR VGND sg13g2_fill_2
XFILLER_43_44 VPWR VGND sg13g2_fill_1
XFILLER_14_959 VPWR VGND sg13g2_decap_8
XFILLER_22_981 VPWR VGND sg13g2_decap_8
X_4952__332 VPWR VGND net332 sg13g2_tiehi
XFILLER_5_679 VPWR VGND sg13g2_decap_8
XFILLER_4_156 VPWR VGND sg13g2_decap_4
XFILLER_1_830 VPWR VGND sg13g2_decap_8
XFILLER_49_812 VPWR VGND sg13g2_decap_8
XFILLER_0_362 VPWR VGND sg13g2_fill_1
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_1_1012 VPWR VGND sg13g2_decap_8
XFILLER_29_591 VPWR VGND sg13g2_decap_8
XFILLER_36_528 VPWR VGND sg13g2_decap_8
XFILLER_16_274 VPWR VGND sg13g2_fill_1
XFILLER_31_211 VPWR VGND sg13g2_decap_4
XFILLER_31_244 VPWR VGND sg13g2_fill_2
X_2820_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\] net758 _0756_ _0488_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_440 VPWR VGND sg13g2_decap_8
XFILLER_9_952 VPWR VGND sg13g2_decap_8
XFILLER_12_491 VPWR VGND sg13g2_fill_2
X_2751_ _0712_ _0714_ _0740_ VPWR VGND sg13g2_nor2_2
XFILLER_31_288 VPWR VGND sg13g2_fill_1
X_2682_ net770 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[2\] _0721_ _0600_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_451 VPWR VGND sg13g2_fill_1
X_4421_ net799 VPWR _2064_ VGND net605 hsync sg13g2_o21ai_1
X_4352_ _1998_ tmds_red.dc_balancing_reg\[2\] _0905_ VPWR VGND sg13g2_nand2_1
X_3303_ _0990_ _0994_ _0995_ VPWR VGND sg13g2_nor2_2
X_4283_ VPWR _1945_ _1944_ VGND sg13g2_inv_1
XFILLER_39_300 VPWR VGND sg13g2_fill_1
X_3234_ _0943_ _0945_ _0946_ _0319_ VPWR VGND sg13g2_nor3_1
XFILLER_39_377 VPWR VGND sg13g2_fill_1
X_3165_ _0894_ _0869_ _0892_ VPWR VGND sg13g2_xnor2_1
X_3096_ net439 green_tmds_par\[2\] net695 serialize.n428\[4\] VPWR VGND sg13g2_mux2_1
XFILLER_22_222 VPWR VGND sg13g2_decap_8
XFILLER_23_745 VPWR VGND sg13g2_fill_1
X_3998_ net612 VPWR _1666_ VGND _1660_ _1665_ sg13g2_o21ai_1
XFILLER_23_778 VPWR VGND sg13g2_fill_2
X_2949_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\] _0790_ _0393_
+ VPWR VGND sg13g2_mux2_1
X_4619_ net665 net717 _0049_ VPWR VGND sg13g2_nor2_1
XFILLER_49_108 VPWR VGND sg13g2_fill_2
XFILLER_38_88 VPWR VGND sg13g2_decap_8
XFILLER_45_314 VPWR VGND sg13g2_fill_1
XFILLER_38_99 VPWR VGND sg13g2_decap_4
XFILLER_18_528 VPWR VGND sg13g2_fill_2
XFILLER_18_539 VPWR VGND sg13g2_decap_8
XFILLER_41_564 VPWR VGND sg13g2_fill_1
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_10_951 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_5_465 VPWR VGND sg13g2_fill_2
XFILLER_49_642 VPWR VGND sg13g2_decap_8
XFILLER_49_631 VPWR VGND sg13g2_fill_2
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_36_347 VPWR VGND sg13g2_fill_2
X_4970_ net305 VGND VPWR _0398_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[1\]
+ _0055_ sg13g2_dfrbpq_1
XFILLER_44_391 VPWR VGND sg13g2_decap_4
X_3921_ _0661_ _1589_ _1590_ VPWR VGND sg13g2_nor2_1
X_3852_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\] net578 _1521_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_575 VPWR VGND sg13g2_decap_8
X_2803_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\] net784 _0752_ _0501_
+ VPWR VGND sg13g2_mux2_1
X_3783_ _1448_ _1449_ _1450_ _1451_ _1452_ VPWR VGND sg13g2_nor4_1
X_2734_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[0\] _0735_ _0562_
+ VPWR VGND sg13g2_mux2_1
X_5170__167 VPWR VGND net167 sg13g2_tiehi
XFILLER_8_292 VPWR VGND sg13g2_decap_8
X_2665_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\] _0713_ _0609_
+ VPWR VGND sg13g2_mux2_1
X_2596_ VPWR _0652_ tmds_green.dc_balancing_reg\[1\] VGND sg13g2_inv_1
X_4404_ VGND VPWR _2022_ _2027_ _2048_ _2026_ sg13g2_a21oi_1
X_4335_ net747 _1989_ _0386_ VPWR VGND sg13g2_nor2_1
X_4266_ VGND VPWR _1928_ _1927_ _1800_ sg13g2_or2_1
X_3217_ _0923_ _0933_ _0307_ VPWR VGND sg13g2_nor2_1
X_4197_ _1859_ _1702_ _1858_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_163 VPWR VGND sg13g2_fill_2
X_3148_ _0877_ tmds_red.n114 _0870_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_859 VPWR VGND sg13g2_fill_2
X_3079_ VGND VPWR serialize.n431\[5\] net697 net413 sg13g2_or2_1
X_4942__342 VPWR VGND net342 sg13g2_tiehi
XFILLER_36_892 VPWR VGND sg13g2_fill_2
XFILLER_35_380 VPWR VGND sg13g2_fill_2
XFILLER_23_553 VPWR VGND sg13g2_fill_1
XFILLER_10_225 VPWR VGND sg13g2_decap_8
XFILLER_6_218 VPWR VGND sg13g2_decap_8
XFILLER_2_413 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_4
XFILLER_3_969 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_fill_2
Xfanout750 net751 net750 VPWR VGND sg13g2_buf_8
XFILLER_46_601 VPWR VGND sg13g2_fill_2
XFILLER_1_28 VPWR VGND sg13g2_decap_4
Xfanout783 ui_in[5] net783 VPWR VGND sg13g2_buf_8
Xfanout761 ui_in[7] net761 VPWR VGND sg13g2_buf_8
Xfanout772 ui_in[6] net772 VPWR VGND sg13g2_buf_8
Xfanout794 ui_in[4] net794 VPWR VGND sg13g2_buf_8
XFILLER_19_837 VPWR VGND sg13g2_fill_1
XFILLER_18_347 VPWR VGND sg13g2_decap_8
XFILLER_34_818 VPWR VGND sg13g2_fill_1
XFILLER_41_394 VPWR VGND sg13g2_fill_1
X_5015__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_6_796 VPWR VGND sg13g2_decap_8
XFILLER_5_273 VPWR VGND sg13g2_fill_2
X_4896__58 VPWR VGND net58 sg13g2_tiehi
X_4120_ _1785_ _1776_ _1777_ VPWR VGND sg13g2_nand2_1
X_4051_ _1714_ VPWR _1716_ VGND _1156_ _1157_ sg13g2_o21ai_1
XFILLER_49_472 VPWR VGND sg13g2_decap_4
X_3002_ _0803_ _0716_ _0744_ VPWR VGND sg13g2_nand2_2
X_4848__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_25_807 VPWR VGND sg13g2_decap_8
XFILLER_36_122 VPWR VGND sg13g2_fill_2
XFILLER_18_870 VPWR VGND sg13g2_decap_4
XFILLER_24_328 VPWR VGND sg13g2_decap_8
X_4953_ net331 VGND VPWR _0381_ tmds_red.n114 net642 sg13g2_dfrbpq_2
X_3904_ _1573_ net594 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\] VPWR
+ VGND sg13g2_nand2b_1
X_4884_ net81 VGND VPWR _0312_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\]
+ _0033_ sg13g2_dfrbpq_1
X_3835_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\] net558 _1504_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_394 VPWR VGND sg13g2_decap_8
X_3766_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[1\] net584 _1435_ VPWR
+ VGND sg13g2_nor2_1
X_2717_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\] net792 _0730_ _0574_
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_15 VPWR VGND sg13g2_fill_1
X_3697_ net615 VPWR _1366_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\]
+ net564 sg13g2_o21ai_1
X_2648_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\] net628 _0701_ VPWR VGND
+ sg13g2_and2_1
X_2579_ VPWR _0635_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[1\] VGND
+ sg13g2_inv_1
X_4318_ _1699_ _1793_ _1399_ _1977_ VPWR VGND sg13g2_nand3_1
X_4249_ VGND VPWR _1904_ _1909_ _1911_ _1907_ sg13g2_a21oi_1
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_19_57 VPWR VGND sg13g2_fill_2
XFILLER_19_79 VPWR VGND sg13g2_fill_2
XFILLER_28_634 VPWR VGND sg13g2_fill_2
X_4862__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_15_306 VPWR VGND sg13g2_decap_8
XFILLER_27_166 VPWR VGND sg13g2_fill_1
XFILLER_23_383 VPWR VGND sg13g2_fill_1
XFILLER_11_534 VPWR VGND sg13g2_decap_4
XFILLER_3_733 VPWR VGND sg13g2_fill_2
Xfanout591 net592 net591 VPWR VGND sg13g2_buf_1
XFILLER_19_612 VPWR VGND sg13g2_decap_8
Xfanout580 net582 net580 VPWR VGND sg13g2_buf_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_19_645 VPWR VGND sg13g2_fill_2
XFILLER_46_475 VPWR VGND sg13g2_fill_1
XFILLER_34_615 VPWR VGND sg13g2_fill_2
XFILLER_30_821 VPWR VGND sg13g2_decap_8
X_3620_ _1288_ _1282_ _1289_ VPWR VGND sg13g2_nor2b_1
X_3551_ _1220_ _1065_ _1218_ VPWR VGND sg13g2_xnor2_1
X_3482_ _1140_ _1119_ _1118_ _1151_ VPWR VGND sg13g2_a21o_1
X_5221_ net804 VGND VPWR serialize.n431\[3\] serialize.n420\[1\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5152_ net312 VGND VPWR _0576_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\]
+ _0224_ sg13g2_dfrbpq_1
X_4877__91 VPWR VGND net91 sg13g2_tiehi
X_4103_ VGND VPWR _1763_ _1765_ _1768_ _1757_ sg13g2_a21oi_1
X_5083_ net367 VGND VPWR _0507_ green_tmds_par\[8\] net637 sg13g2_dfrbpq_1
X_4034_ VPWR _1700_ _1699_ VGND sg13g2_inv_1
XFILLER_37_475 VPWR VGND sg13g2_fill_1
XFILLER_24_125 VPWR VGND sg13g2_fill_2
XFILLER_40_607 VPWR VGND sg13g2_decap_4
X_4936_ net350 VGND VPWR _0364_ videogen.fancy_shader.video_y\[8\] net632 sg13g2_dfrbpq_2
X_4867_ net105 VGND VPWR _0295_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\]
+ _0026_ sg13g2_dfrbpq_1
XFILLER_21_865 VPWR VGND sg13g2_decap_8
X_3818_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\] net588 _1487_ VPWR
+ VGND sg13g2_nor2_1
X_4798_ net691 net742 _0228_ VPWR VGND sg13g2_nor2_1
XFILLER_21_25 VPWR VGND sg13g2_fill_1
X_3749_ _1418_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_0_747 VPWR VGND sg13g2_decap_8
XFILLER_47_206 VPWR VGND sg13g2_decap_4
X_4883__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_46_88 VPWR VGND sg13g2_fill_1
XFILLER_44_957 VPWR VGND sg13g2_decap_8
XFILLER_12_854 VPWR VGND sg13g2_decap_8
XFILLER_8_836 VPWR VGND sg13g2_decap_8
XFILLER_7_324 VPWR VGND sg13g2_fill_2
XFILLER_12_876 VPWR VGND sg13g2_fill_2
XFILLER_12_898 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_fill_2
XFILLER_7_379 VPWR VGND sg13g2_decap_8
X_4874__94 VPWR VGND net94 sg13g2_tiehi
X_4845__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_35_924 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_fill_2
XFILLER_22_607 VPWR VGND sg13g2_fill_1
XFILLER_43_990 VPWR VGND sg13g2_decap_8
X_2982_ _0799_ _0699_ _0722_ VPWR VGND sg13g2_nand2_2
X_4721_ net655 net707 _0151_ VPWR VGND sg13g2_nor2_1
XFILLER_21_128 VPWR VGND sg13g2_decap_8
X_4652_ net669 net722 _0082_ VPWR VGND sg13g2_nor2_1
X_3603_ _1271_ VPWR _1272_ VGND _1263_ _1267_ sg13g2_o21ai_1
X_4583_ net665 net717 _0013_ VPWR VGND sg13g2_nor2_1
X_3534_ _1170_ _1177_ _1202_ _1203_ VPWR VGND sg13g2_or3_1
XFILLER_6_390 VPWR VGND sg13g2_fill_1
X_3465_ _1134_ _1130_ _1131_ _1113_ _1112_ VPWR VGND sg13g2_a22oi_1
X_5204_ net316 VGND VPWR _0628_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\]
+ _0258_ sg13g2_dfrbpq_1
X_3396_ _1065_ _0994_ _1012_ VPWR VGND sg13g2_xnor2_1
X_5135_ net128 VGND VPWR _0559_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[1\]
+ _0207_ sg13g2_dfrbpq_1
X_5066_ net264 VGND VPWR _0003_ videogen.test_lut_thingy.pixel_feeder_inst.state\[1\]
+ net635 sg13g2_dfrbpq_1
X_4017_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\] net556 _1685_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_26_902 VPWR VGND sg13g2_decap_8
XFILLER_26_979 VPWR VGND sg13g2_decap_8
X_4919_ net384 VGND VPWR _0347_ videogen.fancy_shader.n646\[1\] net647 sg13g2_dfrbpq_2
XFILLER_0_522 VPWR VGND sg13g2_decap_8
XFILLER_48_559 VPWR VGND sg13g2_decap_8
X_5122__201 VPWR VGND net201 sg13g2_tiehi
XFILLER_17_968 VPWR VGND sg13g2_decap_8
X_4871__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_28_294 VPWR VGND sg13g2_decap_8
XFILLER_31_448 VPWR VGND sg13g2_fill_2
XFILLER_8_600 VPWR VGND sg13g2_fill_2
X_5092__322 VPWR VGND net322 sg13g2_tiehi
XFILLER_8_633 VPWR VGND sg13g2_fill_2
XFILLER_7_121 VPWR VGND sg13g2_decap_8
X_2612__1 VPWR net405 clknet_1_0__leaf_clk VGND sg13g2_inv_1
XFILLER_7_154 VPWR VGND sg13g2_fill_2
XFILLER_4_883 VPWR VGND sg13g2_decap_8
X_3250_ _0808_ VPWR _0958_ VGND _0647_ _0956_ sg13g2_o21ai_1
XFILLER_26_1000 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_fill_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
X_3181_ _0910_ _0908_ _0909_ _0901_ tmds_red.dc_balancing_reg\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_23_916 VPWR VGND sg13g2_decap_8
X_4997__249 VPWR VGND net249 sg13g2_tiehi
X_5023__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_34_253 VPWR VGND sg13g2_decap_8
XFILLER_34_264 VPWR VGND sg13g2_fill_2
XFILLER_34_275 VPWR VGND sg13g2_decap_8
XFILLER_35_787 VPWR VGND sg13g2_decap_8
XFILLER_22_448 VPWR VGND sg13g2_fill_2
X_4704_ net649 net701 _0134_ VPWR VGND sg13g2_nor2_1
X_2965_ _0794_ _0732_ VPWR VGND _0728_ sg13g2_nand2b_2
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
X_2896_ _0726_ _0772_ _0777_ VPWR VGND sg13g2_nor2_2
X_4635_ net665 net717 _0065_ VPWR VGND sg13g2_nor2_1
XFILLER_8_92 VPWR VGND sg13g2_fill_2
XFILLER_8_81 VPWR VGND sg13g2_fill_1
X_4566_ _2179_ VPWR _2194_ VGND _2176_ _2180_ sg13g2_o21ai_1
X_3517_ VGND VPWR _1185_ _1186_ _1175_ net544 sg13g2_a21oi_2
X_4497_ _2130_ _2127_ _2129_ VPWR VGND sg13g2_xnor2_1
X_4969__307 VPWR VGND net307 sg13g2_tiehi
X_3448_ VGND VPWR _0998_ _1079_ _1117_ _1078_ sg13g2_a21oi_1
X_3379_ videogen.test_lut_thingy.gol_counter_reg\[0\] net746 _0366_ VPWR VGND sg13g2_nor2_1
X_5118_ net217 VGND VPWR _0542_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\]
+ _0190_ sg13g2_dfrbpq_1
X_5049_ net122 VGND VPWR _0477_ videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\]
+ _0134_ sg13g2_dfrbpq_1
XFILLER_26_710 VPWR VGND sg13g2_decap_8
X_4980__286 VPWR VGND net286 sg13g2_tiehi
XFILLER_14_938 VPWR VGND sg13g2_decap_8
XFILLER_25_297 VPWR VGND sg13g2_fill_1
XFILLER_22_960 VPWR VGND sg13g2_decap_8
X_5176__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_5_614 VPWR VGND sg13g2_decap_8
XFILLER_49_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_886 VPWR VGND sg13g2_decap_8
XFILLER_49_868 VPWR VGND sg13g2_decap_8
XFILLER_32_713 VPWR VGND sg13g2_fill_1
XFILLER_9_931 VPWR VGND sg13g2_decap_8
XFILLER_13_982 VPWR VGND sg13g2_decap_8
X_2750_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\] net791 _0739_ _0550_
+ VPWR VGND sg13g2_mux2_1
X_2681_ net760 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[3\] _0721_ _0601_
+ VPWR VGND sg13g2_mux2_1
X_4420_ _2063_ _2062_ VPWR VGND _2057_ sg13g2_nand2b_2
XFILLER_8_474 VPWR VGND sg13g2_fill_2
X_4351_ net571 _1997_ _0510_ VPWR VGND sg13g2_nor2_1
X_3302_ _0994_ _0991_ _0993_ VPWR VGND sg13g2_xnor2_1
X_4282_ _1944_ _1059_ _1858_ VPWR VGND sg13g2_xnor2_1
X_3233_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0941_ _0946_ VPWR VGND
+ sg13g2_and2_1
XFILLER_39_323 VPWR VGND sg13g2_fill_2
XFILLER_39_356 VPWR VGND sg13g2_decap_8
X_3164_ VPWR _0893_ _0892_ VGND sg13g2_inv_1
X_3095_ _0850_ VPWR serialize.n428\[3\] VGND _0669_ net698 sg13g2_o21ai_1
XFILLER_39_389 VPWR VGND sg13g2_fill_2
X_3997_ net615 VPWR _1665_ VGND _1661_ _1664_ sg13g2_o21ai_1
XFILLER_13_37 VPWR VGND sg13g2_decap_8
X_2948_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\] _0790_ _0394_
+ VPWR VGND sg13g2_mux2_1
X_2879_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[1\] _0773_ _0446_
+ VPWR VGND sg13g2_mux2_1
X_4618_ net663 net715 _0048_ VPWR VGND sg13g2_nor2_1
X_4549_ _2178_ _2141_ _2177_ VPWR VGND sg13g2_nand2_1
XFILLER_38_67 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_fill_2
XFILLER_39_890 VPWR VGND sg13g2_fill_2
XFILLER_14_713 VPWR VGND sg13g2_decap_8
XFILLER_41_532 VPWR VGND sg13g2_fill_2
XFILLER_14_757 VPWR VGND sg13g2_decap_4
XFILLER_26_595 VPWR VGND sg13g2_decap_4
XFILLER_10_930 VPWR VGND sg13g2_decap_8
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_23_1014 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_fill_1
XFILLER_17_573 VPWR VGND sg13g2_fill_1
X_3920_ net610 _1565_ _1588_ _1589_ VPWR VGND sg13g2_nor3_1
XFILLER_45_893 VPWR VGND sg13g2_decap_8
X_3851_ net596 VPWR _1520_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\]
+ net566 sg13g2_o21ai_1
X_3782_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\] net554 _1451_ VPWR
+ VGND sg13g2_nor2_1
X_2802_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\] net773 _0752_ _0502_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_727 VPWR VGND sg13g2_fill_1
X_2733_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\] _0735_ _0563_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_271 VPWR VGND sg13g2_decap_8
XFILLER_9_794 VPWR VGND sg13g2_decap_8
X_2664_ _0713_ _0699_ _0711_ VPWR VGND sg13g2_nand2_2
X_2595_ _0651_ net629 VPWR VGND sg13g2_inv_2
X_4403_ _0910_ _2036_ _2041_ _2047_ VPWR VGND sg13g2_nor3_1
X_4334_ VGND VPWR _0906_ _1986_ _1989_ _1988_ sg13g2_a21oi_1
X_4265_ _1927_ _0994_ _1059_ VPWR VGND sg13g2_xnor2_1
X_3216_ _0933_ videogen.fancy_shader.video_x\[8\] _0930_ VPWR VGND sg13g2_xnor2_1
X_4196_ _1005_ _1060_ _1010_ _1858_ VPWR VGND sg13g2_mux2_1
X_3147_ _0663_ _0873_ _0875_ _0876_ VPWR VGND sg13g2_nor3_1
X_3078_ net697 net413 serialize.n431\[4\] VPWR VGND sg13g2_nor2b_1
XFILLER_43_819 VPWR VGND sg13g2_fill_1
XFILLER_23_510 VPWR VGND sg13g2_fill_1
XFILLER_24_36 VPWR VGND sg13g2_decap_8
XFILLER_46_1014 VPWR VGND sg13g2_decap_8
XFILLER_3_948 VPWR VGND sg13g2_decap_8
XFILLER_49_77 VPWR VGND sg13g2_decap_8
Xfanout740 net743 net740 VPWR VGND sg13g2_buf_8
Xfanout751 _0658_ net751 VPWR VGND sg13g2_buf_8
Xfanout784 net785 net784 VPWR VGND sg13g2_buf_8
Xfanout773 net774 net773 VPWR VGND sg13g2_buf_8
Xfanout762 net766 net762 VPWR VGND sg13g2_buf_8
XFILLER_18_304 VPWR VGND sg13g2_decap_8
Xfanout795 net796 net795 VPWR VGND sg13g2_buf_8
X_5043__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_45_167 VPWR VGND sg13g2_fill_2
XFILLER_45_156 VPWR VGND sg13g2_decap_8
XFILLER_27_860 VPWR VGND sg13g2_decap_8
XFILLER_27_871 VPWR VGND sg13g2_fill_2
X_5158__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_14_543 VPWR VGND sg13g2_fill_2
XFILLER_42_885 VPWR VGND sg13g2_decap_8
XFILLER_14_91 VPWR VGND sg13g2_fill_1
XFILLER_2_992 VPWR VGND sg13g2_decap_8
XFILLER_49_451 VPWR VGND sg13g2_decap_8
X_4050_ _1156_ _1157_ _1714_ _1715_ VPWR VGND sg13g2_or3_1
X_3001_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\] _0802_ _0279_
+ VPWR VGND sg13g2_mux2_1
XFILLER_24_307 VPWR VGND sg13g2_decap_8
X_4952_ net332 VGND VPWR _0380_ tmds_red.n100 net642 sg13g2_dfrbpq_2
X_4883_ net83 VGND VPWR _0311_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\]
+ _0032_ sg13g2_dfrbpq_1
X_3903_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\] net559 _1572_ VPWR
+ VGND sg13g2_nor2_1
X_3834_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\] net590 _1503_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_373 VPWR VGND sg13g2_decap_8
X_3765_ net618 VPWR _1434_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[1\]
+ net562 sg13g2_o21ai_1
X_2716_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\] net782 _0730_ _0575_
+ VPWR VGND sg13g2_mux2_1
X_3696_ _1361_ _1362_ _1363_ _1364_ _1365_ VPWR VGND sg13g2_nor4_1
XFILLER_9_591 VPWR VGND sg13g2_decap_4
XFILLER_10_27 VPWR VGND sg13g2_decap_8
X_2647_ _0700_ net545 VPWR VGND _0698_ sg13g2_nand2b_2
XFILLER_10_49 VPWR VGND sg13g2_decap_4
XFILLER_10_38 VPWR VGND sg13g2_fill_1
XFILLER_0_929 VPWR VGND sg13g2_decap_8
X_2578_ VPWR _0634_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[2\] VGND
+ sg13g2_inv_1
X_4317_ _1798_ VPWR _0380_ VGND net747 _1976_ sg13g2_o21ai_1
X_4248_ VGND VPWR _1909_ _1910_ _1907_ _1904_ sg13g2_a21oi_2
X_4179_ _1820_ VPWR _1841_ VGND _1821_ _1826_ sg13g2_o21ai_1
XFILLER_11_524 VPWR VGND sg13g2_decap_4
XFILLER_24_885 VPWR VGND sg13g2_decap_8
XFILLER_11_568 VPWR VGND sg13g2_decap_8
XFILLER_11_579 VPWR VGND sg13g2_fill_1
XFILLER_13_1024 VPWR VGND sg13g2_decap_4
XFILLER_2_266 VPWR VGND sg13g2_decap_8
Xfanout570 _1303_ net570 VPWR VGND sg13g2_buf_8
XFILLER_19_624 VPWR VGND sg13g2_decap_8
Xfanout592 _0687_ net592 VPWR VGND sg13g2_buf_8
Xfanout581 net582 net581 VPWR VGND sg13g2_buf_8
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_46_443 VPWR VGND sg13g2_fill_2
XFILLER_18_123 VPWR VGND sg13g2_fill_1
XFILLER_18_167 VPWR VGND sg13g2_fill_1
XFILLER_46_487 VPWR VGND sg13g2_decap_8
XFILLER_33_104 VPWR VGND sg13g2_decap_8
X_3550_ _1065_ _1218_ _1219_ VPWR VGND sg13g2_nor2_1
X_5220_ net805 VGND VPWR serialize.n431\[2\] serialize.n420\[0\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_6_594 VPWR VGND sg13g2_fill_2
X_3481_ _1119_ _1140_ _1118_ _1150_ VPWR VGND sg13g2_nand3_1
X_5151_ net320 VGND VPWR _0575_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[1\]
+ _0223_ sg13g2_dfrbpq_1
X_5082_ net369 VGND VPWR _0506_ green_tmds_par\[6\] net643 sg13g2_dfrbpq_1
X_4102_ _1763_ _1766_ _1767_ VPWR VGND sg13g2_and2_1
X_4033_ _1699_ _1693_ _1495_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_498 VPWR VGND sg13g2_fill_2
X_4935_ net352 VGND VPWR _0363_ videogen.fancy_shader.video_y\[7\] net632 sg13g2_dfrbpq_2
XFILLER_33_671 VPWR VGND sg13g2_decap_8
X_4866_ net107 VGND VPWR _0294_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[3\]
+ _0025_ sg13g2_dfrbpq_1
XFILLER_32_181 VPWR VGND sg13g2_decap_8
X_4797_ net692 net742 _0227_ VPWR VGND sg13g2_nor2_1
X_3817_ _1486_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_20_365 VPWR VGND sg13g2_fill_1
XFILLER_20_376 VPWR VGND sg13g2_decap_4
XFILLER_21_37 VPWR VGND sg13g2_decap_8
X_3748_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\] net587 _1417_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_21_48 VPWR VGND sg13g2_fill_1
X_3679_ net610 _1347_ _1348_ VPWR VGND sg13g2_nor2_1
X_5033__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_0_726 VPWR VGND sg13g2_decap_8
XFILLER_29_944 VPWR VGND sg13g2_decap_8
XFILLER_28_443 VPWR VGND sg13g2_fill_1
XFILLER_28_465 VPWR VGND sg13g2_fill_1
XFILLER_44_936 VPWR VGND sg13g2_decap_8
XFILLER_43_435 VPWR VGND sg13g2_fill_1
XFILLER_16_627 VPWR VGND sg13g2_decap_8
XFILLER_31_608 VPWR VGND sg13g2_decap_4
XFILLER_43_479 VPWR VGND sg13g2_fill_2
XFILLER_23_192 VPWR VGND sg13g2_decap_4
XFILLER_8_815 VPWR VGND sg13g2_fill_1
XFILLER_7_314 VPWR VGND sg13g2_decap_4
XFILLER_7_336 VPWR VGND sg13g2_fill_2
XFILLER_30_9 VPWR VGND sg13g2_decap_8
XFILLER_39_708 VPWR VGND sg13g2_fill_1
XFILLER_19_410 VPWR VGND sg13g2_fill_1
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_fill_2
XFILLER_34_435 VPWR VGND sg13g2_fill_1
XFILLER_35_969 VPWR VGND sg13g2_decap_8
X_2981_ net787 videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\] _0796_ _0295_
+ VPWR VGND sg13g2_mux2_1
X_4720_ net655 net707 _0150_ VPWR VGND sg13g2_nor2_1
XFILLER_14_181 VPWR VGND sg13g2_fill_2
X_4651_ net670 net721 _0081_ VPWR VGND sg13g2_nor2_1
X_3602_ _1271_ _1269_ _1270_ VPWR VGND sg13g2_xnor2_1
X_4582_ net665 net717 _0012_ VPWR VGND sg13g2_nor2_1
XFILLER_7_892 VPWR VGND sg13g2_decap_8
X_3533_ VPWR VGND _1186_ _1178_ _1184_ _1074_ _1202_ _1075_ sg13g2_a221oi_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_3464_ _1127_ _1128_ _1115_ _1133_ VPWR VGND sg13g2_nand3_1
X_5203_ net373 VGND VPWR _0627_ tmds_blue.dc_balancing_reg\[4\] net638 sg13g2_dfrbpq_2
X_3395_ VPWR _1064_ _1063_ VGND sg13g2_inv_1
X_5134_ net136 VGND VPWR _0558_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[0\]
+ _0206_ sg13g2_dfrbpq_1
XFILLER_29_207 VPWR VGND sg13g2_fill_1
XFILLER_29_218 VPWR VGND sg13g2_fill_2
X_5065_ net263 VGND VPWR _0002_ videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ net635 sg13g2_dfrbpq_1
X_4016_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[0\] net567 _1684_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_26_958 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_decap_8
XFILLER_25_468 VPWR VGND sg13g2_decap_8
XFILLER_40_438 VPWR VGND sg13g2_fill_2
X_4918_ net386 VGND VPWR _0346_ videogen.fancy_shader.n646\[0\] net647 sg13g2_dfrbpq_2
X_4849_ net139 VGND VPWR _0277_ red_tmds_par\[5\] net641 sg13g2_dfrbpq_1
X_4915__392 VPWR VGND net392 sg13g2_tiehi
XFILLER_0_501 VPWR VGND sg13g2_decap_8
X_5085__363 VPWR VGND net363 sg13g2_tiehi
XFILLER_48_538 VPWR VGND sg13g2_decap_8
XFILLER_44_722 VPWR VGND sg13g2_decap_8
XFILLER_17_947 VPWR VGND sg13g2_decap_8
XFILLER_28_273 VPWR VGND sg13g2_fill_2
XFILLER_16_435 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_fill_2
XFILLER_25_991 VPWR VGND sg13g2_decap_8
XFILLER_8_645 VPWR VGND sg13g2_decap_4
XFILLER_11_195 VPWR VGND sg13g2_decap_4
XFILLER_4_862 VPWR VGND sg13g2_decap_8
XFILLER_3_372 VPWR VGND sg13g2_fill_2
X_3180_ tmds_red.dc_balancing_reg\[4\] _0866_ _0909_ VPWR VGND sg13g2_nor2_1
XFILLER_39_538 VPWR VGND sg13g2_fill_2
XFILLER_14_4 VPWR VGND sg13g2_decap_4
XFILLER_47_582 VPWR VGND sg13g2_decap_8
XFILLER_47_571 VPWR VGND sg13g2_decap_4
XFILLER_34_232 VPWR VGND sg13g2_fill_1
XFILLER_35_766 VPWR VGND sg13g2_fill_1
XFILLER_16_980 VPWR VGND sg13g2_decap_8
X_2964_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\] net785 _0793_ _0338_
+ VPWR VGND sg13g2_mux2_1
X_4703_ net679 net731 _0133_ VPWR VGND sg13g2_nor2_1
X_2895_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\] net791 _0776_ _0433_
+ VPWR VGND sg13g2_mux2_1
X_4634_ net665 net717 _0064_ VPWR VGND sg13g2_nor2_1
X_4565_ net572 _2193_ _0626_ VPWR VGND sg13g2_nor2_1
X_3516_ _1172_ _1174_ _1185_ VPWR VGND sg13g2_nor2b_1
X_4496_ _2129_ tmds_green.dc_balancing_reg\[4\] _2128_ VPWR VGND sg13g2_xnor2_1
X_3447_ _0999_ _1000_ _1007_ _1080_ _1116_ VPWR VGND sg13g2_nor4_1
X_3378_ _1038_ _1052_ _0365_ VPWR VGND sg13g2_nor2_1
X_5117_ net221 VGND VPWR _0541_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\]
+ _0189_ sg13g2_dfrbpq_1
X_5048_ net126 VGND VPWR _0476_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\]
+ _0133_ sg13g2_dfrbpq_1
XFILLER_27_36 VPWR VGND sg13g2_fill_1
X_5002__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_14_917 VPWR VGND sg13g2_decap_8
XFILLER_9_409 VPWR VGND sg13g2_decap_8
XFILLER_49_1001 VPWR VGND sg13g2_decap_8
XFILLER_5_659 VPWR VGND sg13g2_decap_8
XFILLER_0_353 VPWR VGND sg13g2_fill_1
XFILLER_1_865 VPWR VGND sg13g2_decap_8
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_0_397 VPWR VGND sg13g2_decap_8
XFILLER_48_346 VPWR VGND sg13g2_decap_8
XFILLER_17_711 VPWR VGND sg13g2_decap_8
XFILLER_17_744 VPWR VGND sg13g2_decap_8
X_4842__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_17_766 VPWR VGND sg13g2_fill_2
XFILLER_32_747 VPWR VGND sg13g2_fill_2
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_13_961 VPWR VGND sg13g2_decap_8
XFILLER_31_246 VPWR VGND sg13g2_fill_1
X_2680_ _0721_ _0720_ VPWR VGND _0719_ sg13g2_nand2b_2
XFILLER_9_987 VPWR VGND sg13g2_decap_8
XFILLER_12_493 VPWR VGND sg13g2_fill_1
X_4350_ _1996_ _0917_ _1997_ VPWR VGND sg13g2_xor2_1
X_3301_ videogen.fancy_shader.n646\[2\] videogen.fancy_shader.video_y\[2\] _0993_
+ VPWR VGND sg13g2_xor2_1
XFILLER_3_180 VPWR VGND sg13g2_fill_2
X_4281_ _1930_ VPWR _1943_ VGND _1937_ _1941_ sg13g2_o21ai_1
X_3232_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] _0941_ _0945_ VPWR VGND
+ sg13g2_nor2_1
X_3163_ _0892_ _0889_ _0891_ VPWR VGND sg13g2_xnor2_1
X_3094_ net436 green_tmds_par\[2\] net696 serialize.n428\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_27_519 VPWR VGND sg13g2_decap_8
XFILLER_35_552 VPWR VGND sg13g2_fill_2
XFILLER_35_574 VPWR VGND sg13g2_fill_2
XFILLER_22_213 VPWR VGND sg13g2_decap_4
XFILLER_23_736 VPWR VGND sg13g2_decap_8
X_3996_ _1663_ VPWR _1664_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\]
+ net554 sg13g2_o21ai_1
X_2947_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\] _0790_ _0395_
+ VPWR VGND sg13g2_mux2_1
X_5075__395 VPWR VGND net395 sg13g2_tiehi
X_2878_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\] _0773_ _0447_
+ VPWR VGND sg13g2_mux2_1
X_4617_ net663 net715 _0047_ VPWR VGND sg13g2_nor2_1
X_4548_ _2166_ VPWR _2177_ VGND _2138_ _2139_ sg13g2_o21ai_1
X_4479_ VPWR _2113_ _2112_ VGND sg13g2_inv_1
XFILLER_18_508 VPWR VGND sg13g2_decap_4
XFILLER_46_839 VPWR VGND sg13g2_decap_8
XFILLER_41_500 VPWR VGND sg13g2_decap_4
XFILLER_14_769 VPWR VGND sg13g2_fill_2
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_10_986 VPWR VGND sg13g2_decap_8
XFILLER_0_172 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_0_183 VPWR VGND sg13g2_fill_2
XFILLER_0_194 VPWR VGND sg13g2_decap_8
XFILLER_48_165 VPWR VGND sg13g2_decap_8
XFILLER_45_872 VPWR VGND sg13g2_decap_8
XFILLER_20_706 VPWR VGND sg13g2_decap_8
X_3850_ VGND VPWR _1519_ _1518_ _1507_ sg13g2_or2_1
X_3781_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\] net564 _1450_ VPWR
+ VGND sg13g2_nor2_1
X_2801_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\] net762 _0752_ _0503_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_739 VPWR VGND sg13g2_fill_2
X_2732_ net767 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\] _0735_ _0564_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
X_2663_ VGND VPWR _0712_ _0710_ net573 sg13g2_or2_1
X_4402_ VGND VPWR _2045_ _2046_ _0512_ net571 sg13g2_a21oi_1
X_2594_ VPWR _0650_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[1\] VGND
+ sg13g2_inv_1
X_4333_ net606 VPWR _1988_ VGND _0906_ _1987_ sg13g2_o21ai_1
X_4264_ VPWR _1926_ _1925_ VGND sg13g2_inv_1
X_3215_ _0932_ videogen.fancy_shader.video_x\[8\] _0930_ VPWR VGND sg13g2_nand2_1
X_4195_ _1855_ _1856_ _1857_ VPWR VGND sg13g2_and2_1
XFILLER_39_165 VPWR VGND sg13g2_fill_1
XFILLER_39_154 VPWR VGND sg13g2_decap_4
X_3146_ _0875_ tmds_red.n100 _0874_ VPWR VGND sg13g2_xnor2_1
X_3077_ net697 net409 serialize.n431\[3\] VPWR VGND sg13g2_nor2b_1
XFILLER_39_187 VPWR VGND sg13g2_decap_4
XFILLER_39_1011 VPWR VGND sg13g2_decap_8
XFILLER_35_382 VPWR VGND sg13g2_fill_1
XFILLER_11_706 VPWR VGND sg13g2_fill_1
XFILLER_23_544 VPWR VGND sg13g2_decap_8
X_3979_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\] net586 _1647_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_3_927 VPWR VGND sg13g2_decap_8
XFILLER_49_56 VPWR VGND sg13g2_decap_8
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
Xfanout730 net732 net730 VPWR VGND sg13g2_buf_8
Xfanout752 net756 net752 VPWR VGND sg13g2_buf_8
Xfanout763 net766 net763 VPWR VGND sg13g2_buf_8
Xfanout774 ui_in[5] net774 VPWR VGND sg13g2_buf_8
Xfanout785 net794 net785 VPWR VGND sg13g2_buf_8
Xfanout796 rst_n net796 VPWR VGND sg13g2_buf_8
XFILLER_41_330 VPWR VGND sg13g2_fill_1
XFILLER_14_577 VPWR VGND sg13g2_decap_8
XFILLER_6_710 VPWR VGND sg13g2_fill_2
XFILLER_10_761 VPWR VGND sg13g2_fill_2
X_5050__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_6_732 VPWR VGND sg13g2_fill_1
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_5_275 VPWR VGND sg13g2_fill_1
XFILLER_2_971 VPWR VGND sg13g2_decap_8
XFILLER_49_485 VPWR VGND sg13g2_fill_1
X_3000_ net776 videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\] _0802_ _0280_
+ VPWR VGND sg13g2_mux2_1
XFILLER_37_614 VPWR VGND sg13g2_fill_2
XFILLER_36_113 VPWR VGND sg13g2_fill_1
XFILLER_36_124 VPWR VGND sg13g2_fill_1
XFILLER_36_135 VPWR VGND sg13g2_fill_2
X_4951_ net333 VGND VPWR _0379_ tmds_red.n102 net641 sg13g2_dfrbpq_2
X_4882_ net85 VGND VPWR _0310_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\]
+ _0031_ sg13g2_dfrbpq_1
X_3902_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\] net581 _1571_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_33_864 VPWR VGND sg13g2_fill_2
X_3833_ net598 VPWR _1502_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\]
+ net576 sg13g2_o21ai_1
XFILLER_32_363 VPWR VGND sg13g2_decap_4
XFILLER_33_886 VPWR VGND sg13g2_decap_8
XFILLER_33_897 VPWR VGND sg13g2_fill_2
XFILLER_20_558 VPWR VGND sg13g2_decap_8
X_3764_ net598 _1427_ _1432_ _1433_ VPWR VGND sg13g2_nor3_1
XFILLER_20_569 VPWR VGND sg13g2_fill_1
X_2715_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[2\] net770 _0730_ _0576_
+ VPWR VGND sg13g2_mux2_1
X_3695_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[2\] net576 _1364_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_581 VPWR VGND sg13g2_decap_4
X_2646_ _0698_ net545 _0699_ VPWR VGND sg13g2_nor2b_2
XFILLER_0_908 VPWR VGND sg13g2_decap_8
X_2577_ VPWR _0633_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[3\] VGND
+ sg13g2_inv_1
X_4895__60 VPWR VGND net60 sg13g2_tiehi
X_4316_ _1799_ VPWR _0379_ VGND net747 _1976_ sg13g2_o21ai_1
X_4247_ VGND VPWR _1890_ _1896_ _1909_ _1908_ sg13g2_a21oi_1
X_4178_ _1840_ _1838_ _1839_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_636 VPWR VGND sg13g2_fill_1
X_3129_ _0859_ tmds_green.n100 _0654_ VPWR VGND sg13g2_nand2_1
XFILLER_27_157 VPWR VGND sg13g2_decap_8
XFILLER_28_669 VPWR VGND sg13g2_fill_1
XFILLER_43_639 VPWR VGND sg13g2_fill_1
XFILLER_43_628 VPWR VGND sg13g2_decap_8
XFILLER_24_831 VPWR VGND sg13g2_decap_4
XFILLER_35_47 VPWR VGND sg13g2_decap_8
XFILLER_23_374 VPWR VGND sg13g2_fill_1
XFILLER_11_547 VPWR VGND sg13g2_fill_2
XFILLER_7_529 VPWR VGND sg13g2_fill_2
XFILLER_13_1003 VPWR VGND sg13g2_decap_8
XFILLER_3_735 VPWR VGND sg13g2_fill_1
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_2_278 VPWR VGND sg13g2_decap_8
Xfanout560 _1300_ net560 VPWR VGND sg13g2_buf_8
Xfanout571 net572 net571 VPWR VGND sg13g2_buf_8
Xfanout593 net594 net593 VPWR VGND sg13g2_buf_8
Xfanout582 _0702_ net582 VPWR VGND sg13g2_buf_8
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_46_422 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_fill_2
XFILLER_19_647 VPWR VGND sg13g2_fill_1
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_19_669 VPWR VGND sg13g2_fill_2
XFILLER_34_606 VPWR VGND sg13g2_fill_1
XFILLER_34_617 VPWR VGND sg13g2_fill_1
X_4925__372 VPWR VGND net372 sg13g2_tiehi
XFILLER_33_127 VPWR VGND sg13g2_fill_2
X_5095__310 VPWR VGND net310 sg13g2_tiehi
XFILLER_15_842 VPWR VGND sg13g2_fill_2
XFILLER_25_80 VPWR VGND sg13g2_fill_2
XFILLER_30_845 VPWR VGND sg13g2_decap_8
XFILLER_30_867 VPWR VGND sg13g2_decap_8
XFILLER_30_878 VPWR VGND sg13g2_fill_1
X_3480_ _1134_ _1136_ _1146_ _1149_ VPWR VGND sg13g2_nor3_1
XFILLER_6_562 VPWR VGND sg13g2_decap_4
XFILLER_44_4 VPWR VGND sg13g2_fill_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_5150_ net351 VGND VPWR _0574_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\]
+ _0222_ sg13g2_dfrbpq_1
X_5081_ net371 VGND VPWR _0505_ green_tmds_par\[2\] net646 sg13g2_dfrbpq_1
X_4101_ _1762_ VPWR _1766_ VGND _1758_ _1765_ sg13g2_o21ai_1
XFILLER_38_923 VPWR VGND sg13g2_fill_1
XFILLER_38_901 VPWR VGND sg13g2_decap_4
X_4032_ VGND VPWR _1299_ _1698_ _0373_ _1596_ sg13g2_a21oi_1
XFILLER_2_73 VPWR VGND sg13g2_fill_2
X_4934_ net354 VGND VPWR _0362_ videogen.fancy_shader.video_y\[6\] net632 sg13g2_dfrbpq_2
XFILLER_24_138 VPWR VGND sg13g2_decap_8
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
XFILLER_21_823 VPWR VGND sg13g2_decap_8
X_4865_ net109 VGND VPWR _0293_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[2\]
+ _0024_ sg13g2_dfrbpq_1
XFILLER_21_834 VPWR VGND sg13g2_fill_1
X_4796_ net690 net742 _0226_ VPWR VGND sg13g2_nor2_1
X_3816_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[1\] net567 _1485_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_399 VPWR VGND sg13g2_fill_1
X_3747_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[1\] net565 _1416_ VPWR
+ VGND sg13g2_nor2_1
X_3678_ net612 _1335_ _1346_ _1347_ VPWR VGND sg13g2_nor3_1
XFILLER_0_705 VPWR VGND sg13g2_decap_8
X_2629_ _0679_ _0680_ _0678_ _0682_ VPWR VGND _0681_ sg13g2_nand4_1
XFILLER_48_709 VPWR VGND sg13g2_fill_1
XFILLER_43_1018 VPWR VGND sg13g2_decap_8
XFILLER_29_923 VPWR VGND sg13g2_decap_8
XFILLER_44_915 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_fill_2
XFILLER_15_116 VPWR VGND sg13g2_fill_2
XFILLER_16_617 VPWR VGND sg13g2_decap_4
XFILLER_16_639 VPWR VGND sg13g2_decap_8
XFILLER_43_447 VPWR VGND sg13g2_decap_8
XFILLER_24_672 VPWR VGND sg13g2_decap_8
XFILLER_24_694 VPWR VGND sg13g2_decap_8
X_4990__267 VPWR VGND net267 sg13g2_tiehi
XFILLER_3_521 VPWR VGND sg13g2_fill_1
XFILLER_3_543 VPWR VGND sg13g2_decap_8
XFILLER_3_576 VPWR VGND sg13g2_decap_8
XFILLER_38_208 VPWR VGND sg13g2_fill_2
XFILLER_4_1023 VPWR VGND sg13g2_decap_4
XFILLER_47_775 VPWR VGND sg13g2_decap_4
XFILLER_47_742 VPWR VGND sg13g2_decap_4
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_35_948 VPWR VGND sg13g2_decap_8
XFILLER_46_296 VPWR VGND sg13g2_fill_1
XFILLER_15_650 VPWR VGND sg13g2_fill_1
X_2980_ VGND VPWR _0650_ _0796_ _0296_ _0798_ sg13g2_a21oi_1
XFILLER_15_683 VPWR VGND sg13g2_decap_8
X_4650_ net670 net721 _0080_ VPWR VGND sg13g2_nor2_1
X_3601_ _1260_ VPWR _1270_ VGND _1250_ _1258_ sg13g2_o21ai_1
X_4581_ net666 net718 _0011_ VPWR VGND sg13g2_nor2_1
X_5200__49 VPWR VGND net49 sg13g2_tiehi
X_3532_ VPWR _1201_ _1200_ VGND sg13g2_inv_1
XFILLER_6_381 VPWR VGND sg13g2_decap_8
X_3463_ _1129_ VPWR _1132_ VGND _1114_ _1126_ sg13g2_o21ai_1
X_5202_ net389 VGND VPWR _0626_ tmds_blue.dc_balancing_reg\[3\] net638 sg13g2_dfrbpq_2
X_5133_ net152 VGND VPWR _0557_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\]
+ _0205_ sg13g2_dfrbpq_1
X_3394_ _1061_ _1062_ _1063_ VPWR VGND sg13g2_and2_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
X_5064_ net262 VGND VPWR _0492_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\]
+ _0149_ sg13g2_dfrbpq_1
X_4015_ _1679_ _1680_ _1681_ _1682_ _1683_ VPWR VGND sg13g2_nor4_1
XFILLER_25_403 VPWR VGND sg13g2_fill_2
XFILLER_26_937 VPWR VGND sg13g2_decap_8
X_4880__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_16_49 VPWR VGND sg13g2_fill_2
XFILLER_25_436 VPWR VGND sg13g2_decap_8
X_4917_ net388 VGND VPWR _0345_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\]
+ _0045_ sg13g2_dfrbpq_1
XFILLER_34_992 VPWR VGND sg13g2_decap_8
X_4848_ net140 VGND VPWR _0276_ red_tmds_par\[3\] net641 sg13g2_dfrbpq_1
XFILLER_5_819 VPWR VGND sg13g2_decap_4
X_4779_ net658 net710 _0209_ VPWR VGND sg13g2_nor2_1
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_557 VPWR VGND sg13g2_decap_8
XFILLER_29_720 VPWR VGND sg13g2_decap_8
XFILLER_28_241 VPWR VGND sg13g2_fill_1
XFILLER_29_764 VPWR VGND sg13g2_decap_4
XFILLER_17_926 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_fill_2
XFILLER_25_970 VPWR VGND sg13g2_decap_8
XFILLER_32_929 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_fill_2
XFILLER_8_602 VPWR VGND sg13g2_fill_1
XFILLER_8_635 VPWR VGND sg13g2_fill_1
XFILLER_11_174 VPWR VGND sg13g2_fill_2
XFILLER_8_668 VPWR VGND sg13g2_decap_4
XFILLER_4_841 VPWR VGND sg13g2_decap_8
XFILLER_3_351 VPWR VGND sg13g2_decap_4
XFILLER_39_517 VPWR VGND sg13g2_decap_8
XFILLER_47_550 VPWR VGND sg13g2_decap_8
XFILLER_19_263 VPWR VGND sg13g2_fill_1
X_2963_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\] net774 _0793_ _0339_
+ VPWR VGND sg13g2_mux2_1
X_4702_ net679 net731 _0132_ VPWR VGND sg13g2_nor2_1
X_2894_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\] net781 _0776_ _0434_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_984 VPWR VGND sg13g2_decap_8
X_4633_ net664 net716 _0063_ VPWR VGND sg13g2_nor2_1
X_4564_ _2183_ _2192_ _2193_ VPWR VGND sg13g2_nor2_1
X_3515_ _1182_ _1181_ _1179_ _1184_ VPWR VGND sg13g2_a21o_1
X_4495_ _2086_ VPWR _2128_ VGND _0653_ _2084_ sg13g2_o21ai_1
X_3446_ _1115_ net609 videogen.fancy_shader.video_x\[8\] VPWR VGND sg13g2_nand2_1
X_3377_ _1052_ videogen.fancy_shader.video_y\[9\] _1051_ VPWR VGND sg13g2_xnor2_1
X_5116_ net225 VGND VPWR _0540_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\]
+ _0188_ sg13g2_dfrbpq_1
X_5047_ net130 VGND VPWR _0475_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\]
+ _0132_ sg13g2_dfrbpq_1
XFILLER_26_756 VPWR VGND sg13g2_decap_4
XFILLER_13_406 VPWR VGND sg13g2_fill_1
XFILLER_26_778 VPWR VGND sg13g2_decap_8
XFILLER_26_789 VPWR VGND sg13g2_fill_2
XFILLER_40_225 VPWR VGND sg13g2_fill_2
XFILLER_43_69 VPWR VGND sg13g2_decap_8
X_4908__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_22_995 VPWR VGND sg13g2_decap_8
XFILLER_1_844 VPWR VGND sg13g2_decap_8
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_0_376 VPWR VGND sg13g2_decap_8
X_5046__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_1_1026 VPWR VGND sg13g2_fill_2
X_4996__251 VPWR VGND net251 sg13g2_tiehi
XFILLER_13_940 VPWR VGND sg13g2_decap_8
XFILLER_40_792 VPWR VGND sg13g2_decap_8
XFILLER_9_966 VPWR VGND sg13g2_decap_8
XFILLER_33_80 VPWR VGND sg13g2_fill_1
X_3300_ videogen.fancy_shader.video_y\[2\] videogen.fancy_shader.n646\[2\] _0992_
+ VPWR VGND sg13g2_and2_1
XFILLER_4_693 VPWR VGND sg13g2_decap_8
X_4280_ _1929_ _1938_ _1928_ _1942_ VPWR VGND _1940_ sg13g2_nand4_1
X_3231_ _0941_ _0943_ _0944_ _0318_ VPWR VGND sg13g2_nor3_1
XFILLER_39_325 VPWR VGND sg13g2_fill_1
X_3162_ _0890_ VPWR _0891_ VGND _0874_ net547 sg13g2_o21ai_1
X_3093_ _0850_ VPWR serialize.n428\[1\] VGND _0668_ net696 sg13g2_o21ai_1
XFILLER_47_380 VPWR VGND sg13g2_fill_1
XFILLER_35_586 VPWR VGND sg13g2_decap_8
XFILLER_22_247 VPWR VGND sg13g2_decap_8
X_3995_ VGND VPWR _0636_ net594 _1663_ _1662_ sg13g2_a21oi_1
X_2946_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\] _0790_ _0396_
+ VPWR VGND sg13g2_mux2_1
X_2877_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\] _0773_ _0448_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_792 VPWR VGND sg13g2_fill_2
X_4616_ net663 net715 _0046_ VPWR VGND sg13g2_nor2_1
X_4547_ _2145_ _2147_ _2176_ VPWR VGND sg13g2_nor2_1
X_4478_ _2087_ _2089_ _2112_ VPWR VGND sg13g2_nor2_1
X_3429_ _1098_ videogen.fancy_shader.video_y\[6\] videogen.fancy_shader.n646\[6\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_38_58 VPWR VGND sg13g2_fill_1
XFILLER_38_47 VPWR VGND sg13g2_decap_4
XFILLER_39_892 VPWR VGND sg13g2_fill_1
XFILLER_41_534 VPWR VGND sg13g2_fill_1
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_9_229 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_5_413 VPWR VGND sg13g2_fill_1
XFILLER_10_965 VPWR VGND sg13g2_decap_8
XFILLER_5_479 VPWR VGND sg13g2_fill_2
XFILLER_48_188 VPWR VGND sg13g2_decap_8
XFILLER_17_542 VPWR VGND sg13g2_decap_8
XFILLER_17_564 VPWR VGND sg13g2_fill_2
XFILLER_17_586 VPWR VGND sg13g2_decap_4
X_3780_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[1\] net576 _1449_ VPWR
+ VGND sg13g2_nor2_1
X_2800_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\] net753 _0752_ _0504_
+ VPWR VGND sg13g2_mux2_1
X_2731_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\] _0735_ _0565_
+ VPWR VGND sg13g2_mux2_1
X_4935__352 VPWR VGND net352 sg13g2_tiehi
X_2662_ net573 _0710_ _0711_ VPWR VGND sg13g2_nor2_2
X_4401_ _2046_ _2035_ _2015_ _2028_ _0913_ VPWR VGND sg13g2_a22oi_1
X_2593_ VPWR _0649_ videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_5_51 VPWR VGND sg13g2_decap_4
X_4332_ _1985_ net547 _1987_ VPWR VGND sg13g2_xor2_1
X_4263_ _1923_ _1924_ _1925_ VPWR VGND sg13g2_and2_1
X_3214_ _0923_ _0930_ _0931_ _0306_ VPWR VGND sg13g2_nor3_1
XFILLER_39_133 VPWR VGND sg13g2_decap_8
X_4194_ VGND VPWR _1856_ _1851_ _1801_ sg13g2_or2_1
X_3145_ tmds_red.n132 tmds_red.n126 _0874_ VPWR VGND sg13g2_xor2_1
X_3076_ net697 net408 serialize.n431\[2\] VPWR VGND sg13g2_nor2b_1
XFILLER_36_851 VPWR VGND sg13g2_decap_8
X_3978_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[0\] net554 _1646_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_23_567 VPWR VGND sg13g2_fill_1
XFILLER_23_578 VPWR VGND sg13g2_decap_4
X_2929_ net765 videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[2\] _0784_ _0407_
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_239 VPWR VGND sg13g2_decap_4
XFILLER_3_906 VPWR VGND sg13g2_decap_8
XFILLER_2_427 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
Xfanout742 net743 net742 VPWR VGND sg13g2_buf_8
Xfanout731 net732 net731 VPWR VGND sg13g2_buf_8
Xfanout720 net723 net720 VPWR VGND sg13g2_buf_8
Xfanout775 net778 net775 VPWR VGND sg13g2_buf_8
Xfanout753 net756 net753 VPWR VGND sg13g2_buf_8
Xfanout764 net766 net764 VPWR VGND sg13g2_buf_8
Xfanout797 net798 net797 VPWR VGND sg13g2_buf_8
Xfanout786 net788 net786 VPWR VGND sg13g2_buf_8
XFILLER_33_309 VPWR VGND sg13g2_fill_2
XFILLER_42_832 VPWR VGND sg13g2_fill_1
XFILLER_27_895 VPWR VGND sg13g2_fill_1
XFILLER_41_320 VPWR VGND sg13g2_decap_4
XFILLER_6_722 VPWR VGND sg13g2_decap_4
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_2_950 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_fill_1
XFILLER_49_497 VPWR VGND sg13g2_decap_4
XFILLER_37_648 VPWR VGND sg13g2_fill_2
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_45_670 VPWR VGND sg13g2_fill_2
XFILLER_17_350 VPWR VGND sg13g2_fill_1
X_4950_ net334 VGND VPWR _0378_ tmds_green.n132 net644 sg13g2_dfrbpq_2
X_3901_ _1566_ _1567_ _1568_ _1569_ _1570_ VPWR VGND sg13g2_nor4_1
X_4881_ net87 VGND VPWR _0309_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\]
+ _0030_ sg13g2_dfrbpq_1
X_3832_ _1497_ _1498_ _1499_ _1500_ _1501_ VPWR VGND sg13g2_nor4_1
XFILLER_20_526 VPWR VGND sg13g2_fill_1
XFILLER_20_537 VPWR VGND sg13g2_decap_8
X_3763_ _1428_ _1429_ _1430_ _1431_ _1432_ VPWR VGND sg13g2_nor4_1
X_2714_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\] net759 _0730_ _0577_
+ VPWR VGND sg13g2_mux2_1
X_3694_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\] net554 _1363_ VPWR
+ VGND sg13g2_nor2_1
X_2645_ _0693_ _0695_ _0685_ _0698_ VPWR VGND sg13g2_nand3_1
X_2576_ VPWR _0632_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[3\] VGND
+ sg13g2_inv_1
X_4315_ net747 _1976_ _0381_ VPWR VGND sg13g2_nor2_1
X_4246_ VGND VPWR _1896_ _1897_ _1908_ _1890_ sg13g2_a21oi_1
XFILLER_19_16 VPWR VGND sg13g2_fill_1
X_4177_ _1839_ _0995_ _1192_ VPWR VGND sg13g2_xnor2_1
X_3128_ net599 net601 _0858_ VPWR VGND sg13g2_xor2_1
X_3059_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0840_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\]
+ _0843_ VPWR VGND sg13g2_nand3_1
X_5057__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_24_810 VPWR VGND sg13g2_decap_8
XFILLER_42_128 VPWR VGND sg13g2_fill_2
XFILLER_24_865 VPWR VGND sg13g2_decap_4
XFILLER_2_202 VPWR VGND sg13g2_fill_2
XFILLER_2_235 VPWR VGND sg13g2_fill_2
Xfanout550 net552 net550 VPWR VGND sg13g2_buf_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
Xfanout572 _0853_ net572 VPWR VGND sg13g2_buf_8
Xfanout561 net565 net561 VPWR VGND sg13g2_buf_8
Xfanout583 _0701_ net583 VPWR VGND sg13g2_buf_8
Xfanout594 _0686_ net594 VPWR VGND sg13g2_buf_8
XFILLER_46_467 VPWR VGND sg13g2_decap_4
XFILLER_46_445 VPWR VGND sg13g2_fill_1
XFILLER_33_139 VPWR VGND sg13g2_fill_2
XFILLER_15_898 VPWR VGND sg13g2_decap_8
XFILLER_30_802 VPWR VGND sg13g2_fill_2
XFILLER_10_581 VPWR VGND sg13g2_fill_1
X_5067__402 VPWR VGND net402 sg13g2_tiehi
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_5080_ net375 VGND VPWR _0504_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\]
+ _0161_ sg13g2_dfrbpq_1
X_4100_ _1750_ _1747_ _1764_ _1765_ VPWR VGND sg13g2_a21o_2
X_4031_ _1398_ _1695_ _1698_ VPWR VGND sg13g2_nor2_1
XFILLER_49_283 VPWR VGND sg13g2_decap_8
XFILLER_38_979 VPWR VGND sg13g2_decap_8
X_4933_ net356 VGND VPWR _0361_ videogen.fancy_shader.video_y\[5\] net632 sg13g2_dfrbpq_2
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
X_4864_ net111 VGND VPWR _0292_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[1\]
+ _0023_ sg13g2_dfrbpq_1
XFILLER_33_695 VPWR VGND sg13g2_decap_4
X_4795_ net690 net742 _0225_ VPWR VGND sg13g2_nor2_1
X_3815_ _1480_ _1481_ _1482_ _1483_ _1484_ VPWR VGND sg13g2_nor4_1
X_3746_ _1411_ _1412_ _1413_ _1414_ _1415_ VPWR VGND sg13g2_nor4_1
X_3677_ net618 _1340_ _1345_ _1346_ VPWR VGND sg13g2_nor3_1
X_2628_ videogen.fancy_shader.video_x\[1\] videogen.fancy_shader.video_x\[0\] _0681_
+ VPWR VGND sg13g2_nor2_1
X_4229_ _1886_ _1888_ _1891_ VPWR VGND _1881_ sg13g2_nand3b_1
XFILLER_46_25 VPWR VGND sg13g2_fill_2
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_28_423 VPWR VGND sg13g2_fill_1
XFILLER_16_607 VPWR VGND sg13g2_fill_2
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_28_478 VPWR VGND sg13g2_decap_8
XFILLER_28_489 VPWR VGND sg13g2_decap_8
XFILLER_24_640 VPWR VGND sg13g2_decap_4
XFILLER_23_183 VPWR VGND sg13g2_fill_1
XFILLER_8_806 VPWR VGND sg13g2_decap_8
XFILLER_7_338 VPWR VGND sg13g2_fill_1
XFILLER_3_555 VPWR VGND sg13g2_decap_8
XFILLER_11_83 VPWR VGND sg13g2_fill_1
XFILLER_4_1002 VPWR VGND sg13g2_decap_8
XFILLER_19_401 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_fill_2
XFILLER_19_445 VPWR VGND sg13g2_decap_4
XFILLER_19_478 VPWR VGND sg13g2_fill_1
XFILLER_35_938 VPWR VGND sg13g2_decap_4
XFILLER_46_286 VPWR VGND sg13g2_decap_4
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_14_183 VPWR VGND sg13g2_fill_1
X_4580_ net665 net717 _0010_ VPWR VGND sg13g2_nor2_1
X_3600_ _1264_ VPWR _1269_ VGND _1250_ _1261_ sg13g2_o21ai_1
X_3531_ _1184_ _1199_ _1200_ VPWR VGND sg13g2_and2_1
X_3462_ _1128_ VPWR _1131_ VGND _1114_ _1126_ sg13g2_o21ai_1
X_3393_ VGND VPWR _1062_ _1060_ _1059_ sg13g2_or2_1
X_5032__180 VPWR VGND net180 sg13g2_tiehi
X_5201_ net33 VGND VPWR _0625_ tmds_blue.dc_balancing_reg\[2\] net639 sg13g2_dfrbpq_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VPWR VGND sg13g2_buf_8
X_5132_ net161 VGND VPWR _0556_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\]
+ _0204_ sg13g2_dfrbpq_1
X_5063_ net55 VGND VPWR _0491_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\]
+ _0148_ sg13g2_dfrbpq_1
X_4014_ net623 VPWR _1682_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[0\]
+ net566 sg13g2_o21ai_1
XFILLER_26_916 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_fill_1
XFILLER_34_971 VPWR VGND sg13g2_decap_8
XFILLER_33_481 VPWR VGND sg13g2_fill_1
X_4916_ net390 VGND VPWR _0344_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\]
+ _0044_ sg13g2_dfrbpq_1
X_5078__383 VPWR VGND net383 sg13g2_tiehi
XFILLER_21_665 VPWR VGND sg13g2_decap_8
XFILLER_33_492 VPWR VGND sg13g2_fill_1
X_4847_ net141 VGND VPWR _0275_ red_tmds_par\[1\] net644 sg13g2_dfrbpq_1
XFILLER_32_49 VPWR VGND sg13g2_fill_1
XFILLER_10_1007 VPWR VGND sg13g2_decap_8
X_4778_ net658 net710 _0208_ VPWR VGND sg13g2_nor2_1
X_3729_ _1398_ _1349_ _1397_ videogen.test_lut_thingy.gol_counter_reg\[2\] _0661_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_536 VPWR VGND sg13g2_decap_8
XFILLER_17_905 VPWR VGND sg13g2_decap_8
XFILLER_44_702 VPWR VGND sg13g2_fill_1
XFILLER_43_201 VPWR VGND sg13g2_decap_4
XFILLER_29_776 VPWR VGND sg13g2_decap_8
XFILLER_29_787 VPWR VGND sg13g2_fill_1
XFILLER_43_256 VPWR VGND sg13g2_decap_4
XFILLER_43_289 VPWR VGND sg13g2_fill_1
XFILLER_12_610 VPWR VGND sg13g2_fill_2
XFILLER_19_1021 VPWR VGND sg13g2_decap_4
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_11_153 VPWR VGND sg13g2_decap_4
XFILLER_11_164 VPWR VGND sg13g2_fill_1
XFILLER_7_135 VPWR VGND sg13g2_decap_8
XFILLER_7_179 VPWR VGND sg13g2_fill_2
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_4_820 VPWR VGND sg13g2_decap_8
XFILLER_4_897 VPWR VGND sg13g2_decap_8
XFILLER_26_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_253 VPWR VGND sg13g2_fill_2
XFILLER_19_286 VPWR VGND sg13g2_fill_2
X_2962_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\] net763 _0793_ _0340_
+ VPWR VGND sg13g2_mux2_1
X_4701_ net680 net730 _0131_ VPWR VGND sg13g2_nor2_1
XFILLER_31_963 VPWR VGND sg13g2_decap_8
X_2893_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\] net771 _0776_ _0435_
+ VPWR VGND sg13g2_mux2_1
X_4632_ net664 net715 _0062_ VPWR VGND sg13g2_nor2_1
XFILLER_30_484 VPWR VGND sg13g2_decap_8
X_4563_ VPWR VGND _2185_ _2057_ _2191_ _2061_ _2192_ _2190_ sg13g2_a221oi_1
X_4494_ VGND VPWR _2101_ _2113_ _2127_ _2126_ sg13g2_a21oi_1
X_3514_ _1181_ _1182_ _1183_ VPWR VGND sg13g2_and2_1
X_3445_ net609 videogen.fancy_shader.video_x\[8\] _1114_ VPWR VGND sg13g2_and2_1
X_3376_ net745 _1050_ _1051_ _0364_ VPWR VGND sg13g2_nor3_1
X_5115_ net229 VGND VPWR _0539_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\]
+ _0187_ sg13g2_dfrbpq_1
XFILLER_38_540 VPWR VGND sg13g2_fill_1
X_5046_ net134 VGND VPWR _0474_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\]
+ _0131_ sg13g2_dfrbpq_1
XFILLER_40_259 VPWR VGND sg13g2_fill_2
XFILLER_22_974 VPWR VGND sg13g2_decap_8
XFILLER_5_606 VPWR VGND sg13g2_decap_4
XFILLER_4_149 VPWR VGND sg13g2_decap_8
XFILLER_0_300 VPWR VGND sg13g2_decap_8
XFILLER_1_823 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_decap_8
XFILLER_1_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_584 VPWR VGND sg13g2_decap_8
XFILLER_44_554 VPWR VGND sg13g2_decap_4
X_5196__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_17_768 VPWR VGND sg13g2_fill_1
XFILLER_17_779 VPWR VGND sg13g2_decap_4
XFILLER_44_587 VPWR VGND sg13g2_decap_4
XFILLER_17_93 VPWR VGND sg13g2_decap_8
XFILLER_31_215 VPWR VGND sg13g2_fill_2
XFILLER_40_760 VPWR VGND sg13g2_fill_2
XFILLER_8_422 VPWR VGND sg13g2_fill_2
XFILLER_8_411 VPWR VGND sg13g2_decap_8
XFILLER_8_400 VPWR VGND sg13g2_decap_8
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_13_996 VPWR VGND sg13g2_decap_8
XFILLER_8_433 VPWR VGND sg13g2_decap_8
X_5053__106 VPWR VGND net106 sg13g2_tiehi
X_5133__152 VPWR VGND net152 sg13g2_tiehi
X_3230_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0940_ _0944_ VPWR VGND
+ sg13g2_nor2_1
X_3161_ _0890_ tmds_red.n126 tmds_red.n132 VPWR VGND sg13g2_nand2b_1
X_3092_ _0850_ green_tmds_par\[1\] net698 VPWR VGND sg13g2_nand2_1
XFILLER_48_893 VPWR VGND sg13g2_decap_8
XFILLER_35_543 VPWR VGND sg13g2_fill_1
XFILLER_35_554 VPWR VGND sg13g2_fill_1
XFILLER_35_565 VPWR VGND sg13g2_decap_4
XFILLER_35_576 VPWR VGND sg13g2_fill_1
X_5001__241 VPWR VGND net241 sg13g2_tiehi
X_3994_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\] net563 _1662_ VPWR
+ VGND sg13g2_nor2_1
X_4858__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_31_771 VPWR VGND sg13g2_fill_1
X_2945_ _0790_ _0781_ VPWR VGND _0728_ sg13g2_nand2b_2
X_2876_ _0773_ _0720_ _0771_ VPWR VGND sg13g2_nand2_2
X_4615_ net689 net739 _0045_ VPWR VGND sg13g2_nor2_1
X_4546_ _2175_ _2171_ _2174_ VPWR VGND sg13g2_xnor2_1
X_4477_ _2109_ _2110_ _2111_ VPWR VGND sg13g2_nor2_1
X_3428_ _1097_ videogen.fancy_shader.video_y\[7\] videogen.fancy_shader.n646\[7\]
+ VPWR VGND sg13g2_xnor2_1
X_3359_ _1040_ _1037_ videogen.fancy_shader.video_y\[3\] _1032_ videogen.fancy_shader.video_y\[2\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_381 VPWR VGND sg13g2_fill_2
X_5029_ net186 VGND VPWR _0457_ videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[0\]
+ _0114_ sg13g2_dfrbpq_1
XFILLER_22_771 VPWR VGND sg13g2_decap_8
XFILLER_10_944 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_370 VPWR VGND sg13g2_fill_2
XFILLER_44_362 VPWR VGND sg13g2_fill_2
XFILLER_32_557 VPWR VGND sg13g2_fill_2
XFILLER_32_568 VPWR VGND sg13g2_decap_8
XFILLER_8_230 VPWR VGND sg13g2_decap_8
X_2730_ _0735_ _0722_ _0732_ VPWR VGND sg13g2_nand2_2
XFILLER_8_263 VPWR VGND sg13g2_decap_4
XFILLER_8_241 VPWR VGND sg13g2_fill_2
X_2661_ _0709_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] _0710_ VPWR VGND
+ _0684_ sg13g2_nand3b_1
XFILLER_8_285 VPWR VGND sg13g2_decap_8
X_4400_ _2043_ _2044_ _0906_ _2045_ VPWR VGND sg13g2_nand3_1
XFILLER_5_30 VPWR VGND sg13g2_decap_8
X_2592_ VPWR _0648_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[1\] VGND sg13g2_inv_1
X_4331_ _1986_ _0910_ _1985_ VPWR VGND sg13g2_xnor2_1
X_4262_ _1873_ _1912_ _1921_ _1924_ VPWR VGND sg13g2_or3_1
X_3213_ net629 _0816_ _0931_ VPWR VGND sg13g2_nor2_1
X_4193_ _1801_ VPWR _1855_ VGND _1851_ _1854_ sg13g2_o21ai_1
X_3144_ _0873_ tmds_red.n114 _0872_ VPWR VGND sg13g2_xnor2_1
X_3075_ net697 net411 serialize.n431\[1\] VPWR VGND sg13g2_nor2b_1
XFILLER_36_885 VPWR VGND sg13g2_decap_8
XFILLER_35_373 VPWR VGND sg13g2_decap_8
X_3977_ net622 VPWR _1645_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\]
+ net576 sg13g2_o21ai_1
XFILLER_11_719 VPWR VGND sg13g2_fill_2
X_2928_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\] _0784_ _0408_
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_218 VPWR VGND sg13g2_decap_8
X_2859_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[2\] _0766_ _0459_
+ VPWR VGND sg13g2_mux2_1
X_4529_ _2060_ _2156_ _2159_ VPWR VGND sg13g2_nor2_1
XFILLER_2_406 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_8 VPWR VGND sg13g2_fill_1
Xfanout721 net723 net721 VPWR VGND sg13g2_buf_8
Xfanout732 net733 net732 VPWR VGND sg13g2_buf_8
Xfanout710 net711 net710 VPWR VGND sg13g2_buf_1
Xfanout754 net755 net754 VPWR VGND sg13g2_buf_8
Xfanout776 net778 net776 VPWR VGND sg13g2_buf_1
Xfanout743 net744 net743 VPWR VGND sg13g2_buf_8
Xfanout765 net766 net765 VPWR VGND sg13g2_buf_8
Xfanout787 net788 net787 VPWR VGND sg13g2_buf_1
XFILLER_19_819 VPWR VGND sg13g2_fill_2
Xfanout798 net806 net798 VPWR VGND sg13g2_buf_2
XFILLER_18_318 VPWR VGND sg13g2_fill_2
XFILLER_27_885 VPWR VGND sg13g2_fill_1
XFILLER_42_899 VPWR VGND sg13g2_decap_4
XFILLER_14_72 VPWR VGND sg13g2_decap_8
XFILLER_5_266 VPWR VGND sg13g2_decap_8
XFILLER_5_299 VPWR VGND sg13g2_decap_4
X_5165__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_49_432 VPWR VGND sg13g2_fill_1
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_fill_1
XFILLER_49_465 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
XFILLER_18_863 VPWR VGND sg13g2_decap_8
XFILLER_33_811 VPWR VGND sg13g2_fill_1
X_3900_ net626 VPWR _1569_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[3\]
+ net559 sg13g2_o21ai_1
X_4880_ net88 VGND VPWR _0308_ videogen.fancy_shader.video_x\[9\] net634 sg13g2_dfrbpq_2
X_3831_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\] net564 _1500_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_33_866 VPWR VGND sg13g2_fill_1
XFILLER_33_877 VPWR VGND sg13g2_fill_2
X_3762_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\] net574 _1431_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_387 VPWR VGND sg13g2_decap_8
XFILLER_13_590 VPWR VGND sg13g2_fill_2
X_2713_ _0707_ _0719_ _0730_ VPWR VGND sg13g2_nor2_2
X_3693_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\] net564 _1362_ VPWR
+ VGND sg13g2_nor2_1
X_2644_ _0697_ _0685_ _0693_ VPWR VGND sg13g2_nand2_1
X_4314_ VGND VPWR _1975_ _1976_ _1971_ _1963_ sg13g2_a21oi_2
X_4245_ _1907_ _1905_ _1906_ VPWR VGND sg13g2_xnor2_1
X_4176_ _1016_ _1013_ _1838_ VPWR VGND sg13g2_xor2_1
XFILLER_19_39 VPWR VGND sg13g2_decap_8
X_3127_ _0857_ net600 tmds_green.n132 VPWR VGND sg13g2_nand2b_1
XFILLER_28_627 VPWR VGND sg13g2_decap_8
X_3058_ VGND VPWR _0835_ _0842_ net16 _0836_ sg13g2_a21oi_1
X_5042__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_35_181 VPWR VGND sg13g2_fill_1
XFILLER_11_516 VPWR VGND sg13g2_decap_4
XFILLER_24_899 VPWR VGND sg13g2_decap_8
XFILLER_3_715 VPWR VGND sg13g2_fill_2
Xfanout551 net552 net551 VPWR VGND sg13g2_buf_1
Xfanout584 net585 net584 VPWR VGND sg13g2_buf_8
Xfanout573 net577 net573 VPWR VGND sg13g2_buf_8
Xfanout562 net565 net562 VPWR VGND sg13g2_buf_1
XFILLER_46_413 VPWR VGND sg13g2_fill_1
Xfanout595 _0659_ net595 VPWR VGND sg13g2_buf_8
XFILLER_18_104 VPWR VGND sg13g2_fill_1
XFILLER_19_638 VPWR VGND sg13g2_decap_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
XFILLER_41_151 VPWR VGND sg13g2_fill_1
XFILLER_25_93 VPWR VGND sg13g2_fill_2
XFILLER_6_520 VPWR VGND sg13g2_decap_4
XFILLER_10_560 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_fill_1
XFILLER_1_280 VPWR VGND sg13g2_fill_2
X_4030_ _1398_ _1495_ _1697_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_75 VPWR VGND sg13g2_fill_1
XFILLER_38_958 VPWR VGND sg13g2_decap_4
XFILLER_17_181 VPWR VGND sg13g2_fill_2
X_4932_ net358 VGND VPWR _0360_ videogen.fancy_shader.video_y\[4\] net633 sg13g2_dfrbpq_2
X_4863_ net113 VGND VPWR _0291_ videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\]
+ _0022_ sg13g2_dfrbpq_1
XFILLER_33_685 VPWR VGND sg13g2_fill_2
X_4794_ net691 net741 _0224_ VPWR VGND sg13g2_nor2_1
X_3814_ net624 VPWR _1483_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\]
+ net578 sg13g2_o21ai_1
XFILLER_21_858 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
X_4976__294 VPWR VGND net294 sg13g2_tiehi
X_3745_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\] net590 _1414_ VPWR
+ VGND sg13g2_nor2_1
X_3676_ _1341_ _1342_ _1343_ _1344_ _1345_ VPWR VGND sg13g2_nor4_1
X_2627_ videogen.fancy_shader.video_x\[8\] videogen.fancy_shader.video_x\[9\] _0680_
+ VPWR VGND sg13g2_nor2b_2
X_4228_ _1881_ _1889_ _1890_ VPWR VGND sg13g2_and2_1
XFILLER_44_906 VPWR VGND sg13g2_fill_1
X_4159_ _1729_ _1018_ _1821_ VPWR VGND sg13g2_xor2_1
XFILLER_29_958 VPWR VGND sg13g2_decap_8
XFILLER_11_313 VPWR VGND sg13g2_fill_2
XFILLER_23_162 VPWR VGND sg13g2_fill_2
XFILLER_11_357 VPWR VGND sg13g2_fill_1
X_4838__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_3_501 VPWR VGND sg13g2_decap_8
X_5049__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_46_221 VPWR VGND sg13g2_fill_2
XFILLER_35_917 VPWR VGND sg13g2_decap_8
XFILLER_43_983 VPWR VGND sg13g2_decap_8
XFILLER_15_696 VPWR VGND sg13g2_decap_4
XFILLER_30_688 VPWR VGND sg13g2_decap_8
X_3530_ _1183_ VPWR _1199_ VGND _1179_ _1186_ sg13g2_o21ai_1
X_3461_ _1127_ _1129_ _1115_ _1130_ VPWR VGND sg13g2_nand3_1
X_3392_ _1061_ _1059_ _1060_ VPWR VGND sg13g2_nand2_1
X_5200_ net49 VGND VPWR _0624_ tmds_blue.dc_balancing_reg\[1\] net639 sg13g2_dfrbpq_2
X_5131_ net165 VGND VPWR _0555_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\]
+ _0203_ sg13g2_dfrbpq_1
X_5062_ net59 VGND VPWR _0490_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\]
+ _0147_ sg13g2_dfrbpq_1
X_4013_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[0\] net579 _1681_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_25_405 VPWR VGND sg13g2_fill_1
XFILLER_34_950 VPWR VGND sg13g2_decap_8
X_4915_ net392 VGND VPWR _0343_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\]
+ _0043_ sg13g2_dfrbpq_1
X_4846_ net142 VGND VPWR _0274_ red_tmds_par\[0\] net644 sg13g2_dfrbpq_1
XFILLER_20_198 VPWR VGND sg13g2_decap_8
X_4777_ net667 net720 _0207_ VPWR VGND sg13g2_nor2_1
XFILLER_4_309 VPWR VGND sg13g2_fill_1
X_3728_ net2 _1396_ _1397_ VPWR VGND sg13g2_and2_1
X_3659_ videogen.test_lut_thingy.pixel_feeder_inst.row\[4\]\[2\] net585 _1328_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_515 VPWR VGND sg13g2_decap_8
X_4868__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_29_711 VPWR VGND sg13g2_decap_4
XFILLER_44_769 VPWR VGND sg13g2_decap_4
XFILLER_43_268 VPWR VGND sg13g2_fill_1
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_12_622 VPWR VGND sg13g2_fill_1
XFILLER_12_633 VPWR VGND sg13g2_fill_1
XFILLER_8_626 VPWR VGND sg13g2_decap_8
XFILLER_7_114 VPWR VGND sg13g2_decap_8
XFILLER_7_103 VPWR VGND sg13g2_fill_2
XFILLER_4_876 VPWR VGND sg13g2_decap_8
XFILLER_47_596 VPWR VGND sg13g2_fill_2
XFILLER_19_298 VPWR VGND sg13g2_decap_4
XFILLER_23_909 VPWR VGND sg13g2_decap_8
X_2961_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\] net752 _0793_ _0341_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_994 VPWR VGND sg13g2_decap_8
X_4700_ net680 net730 _0130_ VPWR VGND sg13g2_nor2_1
XFILLER_31_942 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
X_2892_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\] net759 _0776_ _0436_
+ VPWR VGND sg13g2_mux2_1
X_4631_ net653 net705 _0061_ VPWR VGND sg13g2_nor2_1
XFILLER_8_74 VPWR VGND sg13g2_decap_8
X_4562_ VGND VPWR _2148_ _2181_ _2191_ _2061_ sg13g2_a21oi_1
X_4493_ VPWR VGND net600 _2097_ _2123_ _2102_ _2126_ _2112_ sg13g2_a221oi_1
X_3513_ _1158_ VPWR _1182_ VGND _1169_ _1180_ sg13g2_o21ai_1
XFILLER_6_191 VPWR VGND sg13g2_decap_8
X_3444_ _1109_ VPWR _1113_ VGND _1091_ _1106_ sg13g2_o21ai_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_3375_ _0638_ _0673_ _1043_ _1051_ VPWR VGND sg13g2_nor3_1
X_5114_ net233 VGND VPWR _0538_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\]
+ _0186_ sg13g2_dfrbpq_1
X_5045_ net146 VGND VPWR _0473_ videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[0\]
+ _0130_ sg13g2_dfrbpq_1
XFILLER_26_703 VPWR VGND sg13g2_fill_2
XFILLER_40_227 VPWR VGND sg13g2_fill_1
XFILLER_22_953 VPWR VGND sg13g2_decap_8
X_4829_ _2064_ _2068_ _0614_ VPWR VGND sg13g2_nor2_1
XFILLER_49_1015 VPWR VGND sg13g2_decap_8
XFILLER_4_139 VPWR VGND sg13g2_fill_2
XFILLER_1_802 VPWR VGND sg13g2_decap_8
XFILLER_0_334 VPWR VGND sg13g2_decap_4
XFILLER_1_879 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_17_758 VPWR VGND sg13g2_fill_2
XFILLER_16_268 VPWR VGND sg13g2_fill_1
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_13_975 VPWR VGND sg13g2_decap_8
XFILLER_12_485 VPWR VGND sg13g2_fill_2
XFILLER_39_316 VPWR VGND sg13g2_decap_8
X_3160_ VGND VPWR _0867_ _0882_ _0889_ _0868_ sg13g2_a21oi_1
X_3091_ net423 green_tmds_par\[0\] net696 serialize.n428\[0\] VPWR VGND sg13g2_mux2_1
XFILLER_39_349 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_4
Xhold1 clockdiv.q2 VPWR VGND net406 sg13g2_dlygate4sd3_1
XFILLER_48_872 VPWR VGND sg13g2_decap_8
XFILLER_35_522 VPWR VGND sg13g2_decap_8
XFILLER_35_533 VPWR VGND sg13g2_fill_2
X_3993_ net621 VPWR _1661_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[0\]
+ net575 sg13g2_o21ai_1
X_2944_ VGND VPWR _0636_ _0786_ _0397_ _0789_ sg13g2_a21oi_1
X_2875_ _0772_ _0770_ VPWR VGND net546 sg13g2_nand2b_2
X_4614_ net688 net734 _0044_ VPWR VGND sg13g2_nor2_1
X_4545_ _2174_ tmds_blue.dc_balancing_reg\[4\] _2173_ VPWR VGND sg13g2_xnor2_1
X_4476_ VGND VPWR _2080_ _2090_ _2110_ _2107_ sg13g2_a21oi_1
X_3427_ videogen.fancy_shader.n646\[7\] videogen.fancy_shader.video_y\[7\] _1096_
+ VPWR VGND sg13g2_xor2_1
X_4912__398 VPWR VGND net398 sg13g2_tiehi
X_3358_ _1038_ _1039_ _0358_ VPWR VGND sg13g2_nor2_1
X_5082__369 VPWR VGND net369 sg13g2_tiehi
X_3289_ _0981_ _0982_ _0346_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_883 VPWR VGND sg13g2_decap_8
X_5028_ net188 VGND VPWR _0456_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[3\]
+ _0113_ sg13g2_dfrbpq_1
XFILLER_14_706 VPWR VGND sg13g2_decap_8
XFILLER_41_569 VPWR VGND sg13g2_fill_2
XFILLER_10_923 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_23_1007 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_fill_2
XFILLER_48_179 VPWR VGND sg13g2_decap_4
XFILLER_45_820 VPWR VGND sg13g2_fill_2
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_decap_4
XFILLER_9_732 VPWR VGND sg13g2_decap_8
XFILLER_8_253 VPWR VGND sg13g2_decap_4
XFILLER_12_282 VPWR VGND sg13g2_decap_8
XFILLER_12_293 VPWR VGND sg13g2_fill_2
X_2660_ _0709_ net619 net593 VPWR VGND sg13g2_xnor2_1
X_2591_ _0647_ net628 VPWR VGND sg13g2_inv_2
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4330_ _1985_ tmds_red.n126 _0882_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_97 VPWR VGND sg13g2_decap_8
X_4261_ _1873_ VPWR _1923_ VGND _1912_ _1922_ sg13g2_o21ai_1
X_3212_ net629 _0816_ _0930_ VPWR VGND sg13g2_and2_1
XFILLER_39_113 VPWR VGND sg13g2_fill_2
XFILLER_39_102 VPWR VGND sg13g2_decap_8
X_4192_ _1847_ _1853_ _1854_ VPWR VGND sg13g2_nor2_1
X_5029__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_27_308 VPWR VGND sg13g2_fill_2
X_3143_ _0870_ _0871_ _0872_ VPWR VGND sg13g2_nor2_1
X_3074_ net697 net410 serialize.n431\[0\] VPWR VGND sg13g2_nor2b_1
XFILLER_39_1025 VPWR VGND sg13g2_decap_4
X_3976_ _1643_ VPWR _1644_ VGND _1607_ _1619_ sg13g2_o21ai_1
X_5153__304 VPWR VGND net304 sg13g2_tiehi
X_2927_ _0784_ _0711_ _0781_ VPWR VGND sg13g2_nand2_2
X_2858_ net757 videogen.test_lut_thingy.pixel_feeder_inst.row\[45\]\[3\] _0766_ _0460_
+ VPWR VGND sg13g2_mux2_1
X_2789_ _0726_ _0745_ _0750_ VPWR VGND sg13g2_nor2_2
X_4528_ _2148_ VPWR _2158_ VGND _2149_ _2157_ sg13g2_o21ai_1
XFILLER_46_1007 VPWR VGND sg13g2_decap_8
Xfanout700 net446 net700 VPWR VGND sg13g2_buf_8
X_4459_ _2094_ _2093_ _2092_ VPWR VGND sg13g2_nand2b_1
Xfanout711 net724 net711 VPWR VGND sg13g2_buf_2
Xfanout733 net744 net733 VPWR VGND sg13g2_buf_8
Xfanout722 net723 net722 VPWR VGND sg13g2_buf_8
X_4986__274 VPWR VGND net274 sg13g2_tiehi
Xfanout766 net772 net766 VPWR VGND sg13g2_buf_8
Xfanout744 clockdiv.q1 net744 VPWR VGND sg13g2_buf_8
Xfanout755 net756 net755 VPWR VGND sg13g2_buf_8
Xfanout799 net806 net799 VPWR VGND sg13g2_buf_8
Xfanout777 net778 net777 VPWR VGND sg13g2_buf_8
Xfanout788 net794 net788 VPWR VGND sg13g2_buf_8
XFILLER_45_149 VPWR VGND sg13g2_decap_8
XFILLER_27_853 VPWR VGND sg13g2_decap_8
XFILLER_14_536 VPWR VGND sg13g2_decap_8
XFILLER_42_867 VPWR VGND sg13g2_decap_4
XFILLER_10_720 VPWR VGND sg13g2_fill_2
XFILLER_10_731 VPWR VGND sg13g2_decap_4
X_4889__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_30_94 VPWR VGND sg13g2_decap_8
XFILLER_2_985 VPWR VGND sg13g2_decap_8
XFILLER_49_411 VPWR VGND sg13g2_decap_8
XFILLER_49_444 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_fill_1
XFILLER_33_823 VPWR VGND sg13g2_fill_1
X_3830_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\] net575 _1499_ VPWR
+ VGND sg13g2_nor2_1
X_3761_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\] net561 _1430_ VPWR
+ VGND sg13g2_nor2_1
X_2712_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\] net792 _0729_ _0578_
+ VPWR VGND sg13g2_mux2_1
X_3692_ net598 VPWR _1361_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\]
+ net586 sg13g2_o21ai_1
XFILLER_9_595 VPWR VGND sg13g2_fill_2
X_2643_ _0696_ _0685_ _0695_ VPWR VGND sg13g2_nand2_1
X_4313_ _1697_ _1974_ _1975_ VPWR VGND sg13g2_nor2b_1
X_4244_ _1906_ _1888_ _1892_ VPWR VGND sg13g2_xnor2_1
X_4175_ _1835_ _1833_ _1830_ _1837_ VPWR VGND sg13g2_a21o_1
X_3126_ _0654_ _0855_ _0856_ VPWR VGND sg13g2_and2_1
XFILLER_27_116 VPWR VGND sg13g2_fill_2
XFILLER_43_609 VPWR VGND sg13g2_decap_4
X_3057_ _0842_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\] _0840_ VPWR VGND
+ sg13g2_xnor2_1
XFILLER_23_300 VPWR VGND sg13g2_decap_4
XFILLER_23_333 VPWR VGND sg13g2_decap_8
XFILLER_35_193 VPWR VGND sg13g2_decap_8
XFILLER_11_528 VPWR VGND sg13g2_fill_1
X_3959_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\] net573 _1627_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_13_1017 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_204 VPWR VGND sg13g2_fill_1
XFILLER_2_259 VPWR VGND sg13g2_decap_8
Xfanout574 net577 net574 VPWR VGND sg13g2_buf_8
Xfanout552 net555 net552 VPWR VGND sg13g2_buf_1
Xfanout563 net564 net563 VPWR VGND sg13g2_buf_8
XFILLER_47_948 VPWR VGND sg13g2_decap_8
Xfanout585 net587 net585 VPWR VGND sg13g2_buf_8
Xfanout596 _0645_ net596 VPWR VGND sg13g2_buf_8
XFILLER_46_436 VPWR VGND sg13g2_decap_8
XFILLER_2_782 VPWR VGND sg13g2_decap_8
XFILLER_49_241 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
X_4892__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_18_694 VPWR VGND sg13g2_fill_2
X_4931_ net360 VGND VPWR _0359_ videogen.fancy_shader.video_y\[3\] net633 sg13g2_dfrbpq_2
XFILLER_33_620 VPWR VGND sg13g2_decap_8
X_4862_ net115 VGND VPWR _0290_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[3\]
+ _0021_ sg13g2_dfrbpq_1
XFILLER_32_141 VPWR VGND sg13g2_fill_2
XFILLER_33_642 VPWR VGND sg13g2_decap_8
XFILLER_33_664 VPWR VGND sg13g2_decap_8
X_3813_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\] net589 _1482_ VPWR
+ VGND sg13g2_nor2_1
X_4793_ net690 net741 _0223_ VPWR VGND sg13g2_nor2_1
XFILLER_20_358 VPWR VGND sg13g2_decap_8
X_3744_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[1\] net568 _1413_ VPWR
+ VGND sg13g2_nor2_1
X_3675_ videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[2\] net550 _1344_ VPWR
+ VGND sg13g2_nor2_1
X_2626_ _0651_ videogen.fancy_shader.video_x\[3\] videogen.fancy_shader.video_x\[2\]
+ _0679_ VPWR VGND sg13g2_nor3_1
XFILLER_0_719 VPWR VGND sg13g2_decap_8
X_4227_ _1886_ _1888_ _1884_ _1889_ VPWR VGND sg13g2_nand3_1
XFILLER_28_403 VPWR VGND sg13g2_fill_2
XFILLER_29_937 VPWR VGND sg13g2_decap_8
X_4158_ VGND VPWR _1820_ _1819_ _1818_ sg13g2_or2_1
XFILLER_28_436 VPWR VGND sg13g2_decap_8
XFILLER_44_929 VPWR VGND sg13g2_decap_8
X_3109_ net431 red_tmds_par\[7\] net696 serialize.n427\[7\] VPWR VGND sg13g2_mux2_1
X_4089_ _1754_ _1705_ _1753_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_428 VPWR VGND sg13g2_decap_8
XFILLER_23_196 VPWR VGND sg13g2_fill_2
XFILLER_7_318 VPWR VGND sg13g2_fill_1
XFILLER_7_307 VPWR VGND sg13g2_decap_8
XFILLER_46_233 VPWR VGND sg13g2_fill_1
XFILLER_19_425 VPWR VGND sg13g2_decap_8
XFILLER_28_992 VPWR VGND sg13g2_decap_8
XFILLER_36_60 VPWR VGND sg13g2_fill_1
XFILLER_43_962 VPWR VGND sg13g2_decap_8
XFILLER_14_163 VPWR VGND sg13g2_fill_1
XFILLER_30_634 VPWR VGND sg13g2_decap_4
XFILLER_30_645 VPWR VGND sg13g2_decap_4
XFILLER_7_885 VPWR VGND sg13g2_decap_8
X_3460_ _1129_ videogen.fancy_shader.n646\[9\] videogen.fancy_shader.video_x\[9\]
+ VPWR VGND sg13g2_xnor2_1
X_3391_ _1005_ _1004_ _1060_ VPWR VGND sg13g2_xor2_1
X_5130_ net169 VGND VPWR _0554_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\]
+ _0202_ sg13g2_dfrbpq_1
X_5061_ net63 VGND VPWR _0489_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\]
+ _0146_ sg13g2_dfrbpq_1
X_4012_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\] net557 _1680_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_25_417 VPWR VGND sg13g2_fill_2
XFILLER_18_491 VPWR VGND sg13g2_decap_4
X_4914_ net394 VGND VPWR _0342_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\]
+ _0042_ sg13g2_dfrbpq_1
X_4845_ net143 VGND VPWR _0273_ green_tmds_par\[7\] net645 sg13g2_dfrbpq_1
XFILLER_21_645 VPWR VGND sg13g2_fill_2
XFILLER_21_689 VPWR VGND sg13g2_decap_4
X_4776_ net668 net719 _0206_ VPWR VGND sg13g2_nor2_1
X_3727_ _1395_ VPWR _1396_ VGND _1360_ _1371_ sg13g2_o21ai_1
X_3658_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\] net574 _1327_ VPWR
+ VGND sg13g2_nor2_1
X_5011__222 VPWR VGND net222 sg13g2_tiehi
X_3589_ VPWR VGND _1256_ _1090_ _1254_ _1148_ _1258_ _1173_ sg13g2_a221oi_1
X_2609_ VPWR _0665_ tmds_red.dc_balancing_reg\[1\] VGND sg13g2_inv_1
XFILLER_28_222 VPWR VGND sg13g2_fill_1
XFILLER_29_734 VPWR VGND sg13g2_fill_1
XFILLER_16_406 VPWR VGND sg13g2_fill_1
XFILLER_16_428 VPWR VGND sg13g2_decap_8
X_4922__378 VPWR VGND net378 sg13g2_tiehi
XFILLER_25_984 VPWR VGND sg13g2_decap_8
XFILLER_40_932 VPWR VGND sg13g2_fill_2
XFILLER_24_483 VPWR VGND sg13g2_fill_2
XFILLER_11_133 VPWR VGND sg13g2_decap_4
XFILLER_12_656 VPWR VGND sg13g2_decap_4
XFILLER_7_148 VPWR VGND sg13g2_fill_2
XFILLER_11_199 VPWR VGND sg13g2_fill_2
XFILLER_22_73 VPWR VGND sg13g2_decap_8
XFILLER_22_84 VPWR VGND sg13g2_decap_4
XFILLER_4_855 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_39_509 VPWR VGND sg13g2_decap_4
X_5166__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_47_531 VPWR VGND sg13g2_fill_1
XFILLER_14_8 VPWR VGND sg13g2_fill_1
XFILLER_47_564 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_47_575 VPWR VGND sg13g2_fill_2
XFILLER_34_247 VPWR VGND sg13g2_fill_2
X_2960_ _0700_ _0726_ _0793_ VPWR VGND sg13g2_nor2_2
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_31_921 VPWR VGND sg13g2_decap_8
XFILLER_42_291 VPWR VGND sg13g2_decap_4
X_2891_ _0737_ _0772_ _0776_ VPWR VGND sg13g2_nor2_2
XFILLER_8_20 VPWR VGND sg13g2_decap_8
X_4630_ net652 net704 _0060_ VPWR VGND sg13g2_nor2_1
XFILLER_30_464 VPWR VGND sg13g2_decap_4
XFILLER_31_998 VPWR VGND sg13g2_decap_8
X_4561_ _2190_ _2189_ _2188_ VPWR VGND sg13g2_nand2b_1
X_4492_ VGND VPWR _2125_ _2124_ _2097_ sg13g2_or2_1
XFILLER_7_682 VPWR VGND sg13g2_decap_4
XFILLER_6_170 VPWR VGND sg13g2_fill_2
X_3512_ _1149_ _1158_ _1180_ _1181_ VPWR VGND sg13g2_or3_1
X_3443_ _1107_ _1108_ _1092_ _1112_ VPWR VGND sg13g2_nand3_1
X_5113_ net236 VGND VPWR _0537_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\]
+ _0185_ sg13g2_dfrbpq_1
X_3374_ videogen.fancy_shader.video_y\[8\] _1049_ _1050_ VPWR VGND sg13g2_nor2_1
XFILLER_33_0 VPWR VGND sg13g2_decap_4
X_5044_ net150 VGND VPWR _0472_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\]
+ _0129_ sg13g2_dfrbpq_1
XFILLER_38_586 VPWR VGND sg13g2_decap_4
XFILLER_25_269 VPWR VGND sg13g2_fill_2
XFILLER_22_932 VPWR VGND sg13g2_decap_8
X_4828_ _2064_ _2068_ _0613_ VPWR VGND sg13g2_nor2_1
X_5039__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_21_464 VPWR VGND sg13g2_fill_1
X_4759_ net683 net734 _0189_ VPWR VGND sg13g2_nor2_1
X_4835__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_1_858 VPWR VGND sg13g2_decap_8
XFILLER_17_704 VPWR VGND sg13g2_decap_8
XFILLER_29_542 VPWR VGND sg13g2_fill_2
XFILLER_17_737 VPWR VGND sg13g2_decap_8
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_13_954 VPWR VGND sg13g2_decap_8
XFILLER_12_442 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_4
XFILLER_4_652 VPWR VGND sg13g2_decap_8
XFILLER_4_663 VPWR VGND sg13g2_fill_1
XFILLER_3_173 VPWR VGND sg13g2_decap_8
X_3090_ blue_tmds_par\[9\] net694 serialize.n429\[9\] VPWR VGND sg13g2_and2_1
XFILLER_0_880 VPWR VGND sg13g2_decap_8
Xhold2 _0623_ VPWR VGND net407 sg13g2_dlygate4sd3_1
XFILLER_48_851 VPWR VGND sg13g2_decap_8
XFILLER_47_394 VPWR VGND sg13g2_decap_4
X_3992_ net621 _1656_ _1657_ _1659_ _1660_ VPWR VGND sg13g2_nor4_1
XFILLER_22_206 VPWR VGND sg13g2_decap_8
XFILLER_22_217 VPWR VGND sg13g2_fill_1
X_2943_ net787 _0786_ _0789_ VPWR VGND sg13g2_nor2_1
XFILLER_31_762 VPWR VGND sg13g2_decap_8
X_2874_ net546 _0770_ _0771_ VPWR VGND sg13g2_nor2b_2
XFILLER_30_261 VPWR VGND sg13g2_fill_1
X_4613_ net689 net740 _0043_ VPWR VGND sg13g2_nor2_1
X_4544_ _2172_ VPWR _2173_ VGND tmds_blue.dc_balancing_reg\[3\] _2140_ sg13g2_o21ai_1
X_4475_ _2109_ _0863_ _2108_ VPWR VGND sg13g2_nand2_1
X_3426_ VGND VPWR _1069_ _1084_ _1095_ _1083_ sg13g2_a21oi_1
X_3357_ _1039_ _0640_ _1033_ VPWR VGND sg13g2_xnor2_1
X_3288_ VGND VPWR _0643_ _0942_ _0982_ net750 sg13g2_a21oi_1
X_5027_ net190 VGND VPWR _0455_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\]
+ _0112_ sg13g2_dfrbpq_1
XFILLER_26_545 VPWR VGND sg13g2_decap_4
XFILLER_41_504 VPWR VGND sg13g2_fill_1
XFILLER_26_567 VPWR VGND sg13g2_fill_1
XFILLER_10_902 VPWR VGND sg13g2_decap_8
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
XFILLER_22_740 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_fill_1
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_10_979 VPWR VGND sg13g2_decap_8
XFILLER_1_611 VPWR VGND sg13g2_fill_1
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_48_125 VPWR VGND sg13g2_decap_8
XFILLER_29_372 VPWR VGND sg13g2_fill_1
XFILLER_45_865 VPWR VGND sg13g2_fill_2
XFILLER_44_82 VPWR VGND sg13g2_fill_1
XFILLER_13_740 VPWR VGND sg13g2_fill_2
XFILLER_32_559 VPWR VGND sg13g2_fill_1
XFILLER_40_581 VPWR VGND sg13g2_decap_8
XFILLER_13_773 VPWR VGND sg13g2_fill_2
XFILLER_13_795 VPWR VGND sg13g2_decap_8
X_2590_ _0646_ net619 VPWR VGND sg13g2_inv_2
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_4260_ _1922_ _1919_ _1920_ _1915_ _1913_ VPWR VGND sg13g2_a22oi_1
X_3211_ _0816_ _0923_ _0929_ _0305_ VPWR VGND sg13g2_nor3_1
X_4191_ _1853_ _1849_ _1852_ VPWR VGND sg13g2_nand2_2
X_3142_ tmds_red.n126 tmds_red.n132 _0871_ VPWR VGND sg13g2_nor2_1
XFILLER_39_158 VPWR VGND sg13g2_fill_1
XFILLER_39_147 VPWR VGND sg13g2_decap_8
X_3073_ net412 net695 serialize.n433\[0\] VPWR VGND sg13g2_nor2_1
XFILLER_36_821 VPWR VGND sg13g2_fill_2
XFILLER_35_320 VPWR VGND sg13g2_decap_4
XFILLER_35_331 VPWR VGND sg13g2_fill_1
XFILLER_39_1004 VPWR VGND sg13g2_decap_8
XFILLER_36_898 VPWR VGND sg13g2_decap_8
XFILLER_36_865 VPWR VGND sg13g2_decap_4
X_3975_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[5\] _1642_ _1643_ VPWR VGND
+ sg13g2_nor2_1
X_2926_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\] _0783_ _0409_
+ VPWR VGND sg13g2_mux2_1
X_2857_ _0766_ _0757_ VPWR VGND _0728_ sg13g2_nand2b_2
XFILLER_31_592 VPWR VGND sg13g2_fill_2
X_2788_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\] net785 _0749_ _0522_
+ VPWR VGND sg13g2_mux2_1
X_4527_ _2134_ net602 _2157_ VPWR VGND sg13g2_nor2b_1
X_4458_ _2093_ _2090_ _2091_ VPWR VGND sg13g2_nand2_1
XFILLER_49_49 VPWR VGND sg13g2_decap_8
Xfanout701 net703 net701 VPWR VGND sg13g2_buf_8
X_3409_ videogen.fancy_shader.n646\[5\] videogen.fancy_shader.video_x\[5\] _1078_
+ VPWR VGND sg13g2_nor2_1
Xfanout712 net714 net712 VPWR VGND sg13g2_buf_8
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_8
Xfanout734 net738 net734 VPWR VGND sg13g2_buf_8
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
Xfanout767 net769 net767 VPWR VGND sg13g2_buf_8
Xfanout756 ui_in[7] net756 VPWR VGND sg13g2_buf_8
X_4389_ _2031_ _2033_ _2034_ VPWR VGND sg13g2_nor2b_1
Xfanout789 net790 net789 VPWR VGND sg13g2_buf_8
Xfanout778 ui_in[5] net778 VPWR VGND sg13g2_buf_8
X_5123__197 VPWR VGND net197 sg13g2_tiehi
X_4993__257 VPWR VGND net257 sg13g2_tiehi
XFILLER_14_96 VPWR VGND sg13g2_decap_4
XFILLER_5_202 VPWR VGND sg13g2_decap_8
XFILLER_6_769 VPWR VGND sg13g2_fill_2
XFILLER_2_964 VPWR VGND sg13g2_decap_8
X_4965__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_36_106 VPWR VGND sg13g2_fill_1
XFILLER_33_802 VPWR VGND sg13g2_decap_8
XFILLER_44_194 VPWR VGND sg13g2_decap_4
XFILLER_32_345 VPWR VGND sg13g2_decap_4
XFILLER_33_857 VPWR VGND sg13g2_decap_8
XFILLER_33_879 VPWR VGND sg13g2_fill_1
X_3760_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\] net584 _1429_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_367 VPWR VGND sg13g2_fill_2
X_2711_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[1\] net782 _0729_ _0579_
+ VPWR VGND sg13g2_mux2_1
X_3691_ net625 _1354_ _1359_ _1360_ VPWR VGND sg13g2_nor3_1
XFILLER_9_585 VPWR VGND sg13g2_fill_2
X_2642_ _0695_ net610 _0692_ VPWR VGND sg13g2_xnor2_1
X_4312_ VGND VPWR _1398_ _1700_ _1974_ _1973_ sg13g2_a21oi_1
X_4243_ _1877_ _1894_ _1898_ _1905_ VPWR VGND sg13g2_nor3_1
X_4174_ _1836_ _1830_ _1833_ VPWR VGND sg13g2_nand2_1
X_3125_ tmds_green.dc_balancing_reg\[0\] tmds_green.dc_balancing_reg\[1\] tmds_green.dc_balancing_reg\[3\]
+ tmds_green.dc_balancing_reg\[2\] _0855_ VPWR VGND sg13g2_nor4_1
X_3056_ VGND VPWR _0835_ _0841_ net15 _0836_ sg13g2_a21oi_1
XFILLER_36_651 VPWR VGND sg13g2_decap_4
XFILLER_24_824 VPWR VGND sg13g2_decap_8
XFILLER_24_835 VPWR VGND sg13g2_fill_2
XFILLER_23_367 VPWR VGND sg13g2_decap_8
X_3958_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\] net561 _1626_ VPWR
+ VGND sg13g2_nor2_1
X_2909_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[1\] net778 _0779_ _0422_
+ VPWR VGND sg13g2_mux2_1
X_3889_ _1554_ _1555_ _1556_ _1557_ _1558_ VPWR VGND sg13g2_nor4_1
XFILLER_3_717 VPWR VGND sg13g2_fill_1
XFILLER_2_216 VPWR VGND sg13g2_decap_4
Xfanout564 net565 net564 VPWR VGND sg13g2_buf_8
Xfanout553 net554 net553 VPWR VGND sg13g2_buf_8
Xfanout575 net576 net575 VPWR VGND sg13g2_buf_8
XFILLER_47_927 VPWR VGND sg13g2_decap_8
Xfanout597 _0645_ net597 VPWR VGND sg13g2_buf_8
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_8
X_5021__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_15_835 VPWR VGND sg13g2_decap_8
XFILLER_26_150 VPWR VGND sg13g2_decap_4
XFILLER_27_673 VPWR VGND sg13g2_decap_4
XFILLER_15_868 VPWR VGND sg13g2_decap_4
XFILLER_25_51 VPWR VGND sg13g2_fill_1
XFILLER_25_62 VPWR VGND sg13g2_fill_1
XFILLER_41_142 VPWR VGND sg13g2_decap_8
XFILLER_25_73 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_fill_1
XFILLER_41_94 VPWR VGND sg13g2_decap_4
X_4932__358 VPWR VGND net358 sg13g2_tiehi
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
X_5169__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_37_7 VPWR VGND sg13g2_fill_1
XFILLER_2_761 VPWR VGND sg13g2_decap_8
XFILLER_49_220 VPWR VGND sg13g2_decap_8
XFILLER_38_905 VPWR VGND sg13g2_fill_1
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_49_275 VPWR VGND sg13g2_decap_4
XFILLER_38_938 VPWR VGND sg13g2_fill_2
XFILLER_2_66 VPWR VGND sg13g2_decap_8
XFILLER_49_297 VPWR VGND sg13g2_fill_1
XFILLER_2_99 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_fill_2
XFILLER_46_993 VPWR VGND sg13g2_decap_8
XFILLER_45_470 VPWR VGND sg13g2_fill_2
X_4930_ net362 VGND VPWR _0358_ videogen.fancy_shader.video_y\[2\] net633 sg13g2_dfrbpq_2
X_4861_ net117 VGND VPWR _0289_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[2\]
+ _0020_ sg13g2_dfrbpq_1
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
XFILLER_17_183 VPWR VGND sg13g2_fill_1
X_3812_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\] net566 _1481_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_304 VPWR VGND sg13g2_fill_2
X_4792_ net691 net741 _0222_ VPWR VGND sg13g2_nor2_1
X_3743_ videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\] net580 _1412_ VPWR
+ VGND sg13g2_nor2_1
X_3674_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\] net575 _1343_ VPWR
+ VGND sg13g2_nor2_1
X_2625_ videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\] videogen.fancy_shader.video_x\[4\]
+ _0678_ VPWR VGND sg13g2_nor3_1
X_4226_ _1888_ _1158_ _1887_ VPWR VGND sg13g2_xnor2_1
X_4157_ VGND VPWR _1810_ _1814_ _1819_ _1804_ sg13g2_a21oi_1
XFILLER_29_916 VPWR VGND sg13g2_decap_8
X_3108_ net430 red_tmds_par\[6\] net695 serialize.n427\[6\] VPWR VGND sg13g2_mux2_1
XFILLER_37_960 VPWR VGND sg13g2_decap_4
X_4088_ VGND VPWR _1747_ _1750_ _1753_ _1752_ sg13g2_a21oi_1
XFILLER_37_993 VPWR VGND sg13g2_decap_8
X_3039_ VGND VPWR net595 net12 _0693_ net549 sg13g2_a21oi_2
XFILLER_12_816 VPWR VGND sg13g2_fill_2
XFILLER_24_665 VPWR VGND sg13g2_decap_8
XFILLER_24_687 VPWR VGND sg13g2_decap_8
XFILLER_11_315 VPWR VGND sg13g2_fill_1
X_5060__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_3_569 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1016 VPWR VGND sg13g2_decap_8
XFILLER_47_746 VPWR VGND sg13g2_fill_2
XFILLER_46_201 VPWR VGND sg13g2_fill_2
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_28_971 VPWR VGND sg13g2_decap_8
XFILLER_43_941 VPWR VGND sg13g2_decap_8
XFILLER_15_676 VPWR VGND sg13g2_decap_8
XFILLER_7_842 VPWR VGND sg13g2_decap_4
XFILLER_10_381 VPWR VGND sg13g2_decap_4
X_3390_ _1059_ _0987_ _0988_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_4 VPWR VGND sg13g2_fill_2
X_5060_ net67 VGND VPWR _0488_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[3\]
+ _0145_ sg13g2_dfrbpq_1
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
X_4011_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\] net589 _1679_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_19_993 VPWR VGND sg13g2_decap_8
X_4913_ net396 VGND VPWR _0341_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\]
+ _0041_ sg13g2_dfrbpq_1
XFILLER_34_985 VPWR VGND sg13g2_decap_8
X_4844_ net144 VGND VPWR _0272_ green_tmds_par\[1\] net643 sg13g2_dfrbpq_1
X_4775_ net657 net709 _0205_ VPWR VGND sg13g2_nor2_1
XFILLER_21_679 VPWR VGND sg13g2_fill_2
X_3726_ _1394_ net610 _1395_ VPWR VGND sg13g2_nor2b_1
X_3657_ videogen.test_lut_thingy.pixel_feeder_inst.row\[5\]\[2\] net562 _1326_ VPWR
+ VGND sg13g2_nor2_1
X_3588_ _1257_ _1254_ _1256_ _1173_ _1148_ VPWR VGND sg13g2_a22oi_1
X_2608_ VPWR _0664_ tmds_red.dc_balancing_reg\[4\] VGND sg13g2_inv_1
X_5189_ net203 VGND VPWR _0613_ blue_tmds_par\[3\] net637 sg13g2_dfrbpq_1
X_4209_ _1869_ _1192_ _1871_ VPWR VGND sg13g2_xor2_1
XFILLER_17_919 VPWR VGND sg13g2_decap_8
XFILLER_28_234 VPWR VGND sg13g2_decap_8
XFILLER_24_451 VPWR VGND sg13g2_fill_1
XFILLER_25_963 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_fill_1
XFILLER_40_999 VPWR VGND sg13g2_decap_8
XFILLER_4_801 VPWR VGND sg13g2_decap_4
XFILLER_4_834 VPWR VGND sg13g2_decap_8
XFILLER_3_344 VPWR VGND sg13g2_fill_2
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_543 VPWR VGND sg13g2_decap_8
XFILLER_47_598 VPWR VGND sg13g2_fill_1
XFILLER_16_952 VPWR VGND sg13g2_decap_8
XFILLER_31_900 VPWR VGND sg13g2_decap_8
X_2890_ net792 videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\] _0775_ _0437_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_473 VPWR VGND sg13g2_fill_1
X_5173__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_31_977 VPWR VGND sg13g2_decap_8
X_4560_ _2156_ _2187_ _2134_ _2189_ VPWR VGND sg13g2_nand3_1
XFILLER_30_498 VPWR VGND sg13g2_fill_1
X_4491_ _2114_ _2123_ net600 _2124_ VPWR VGND sg13g2_nand3_1
X_3511_ net544 _1170_ _1176_ _1180_ VPWR VGND sg13g2_nor3_1
X_3442_ _1108_ VPWR _1111_ VGND _1091_ _1106_ sg13g2_o21ai_1
XFILLER_40_2 VPWR VGND sg13g2_fill_1
X_3373_ net745 _1048_ _1049_ _0363_ VPWR VGND sg13g2_nor3_1
X_5112_ net240 VGND VPWR _0536_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\]
+ _0184_ sg13g2_dfrbpq_1
X_5043_ net157 VGND VPWR _0471_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[2\]
+ _0128_ sg13g2_dfrbpq_1
XFILLER_25_237 VPWR VGND sg13g2_decap_4
XFILLER_26_749 VPWR VGND sg13g2_decap_8
XFILLER_22_911 VPWR VGND sg13g2_decap_8
XFILLER_40_218 VPWR VGND sg13g2_fill_2
X_4827_ net657 net709 _0257_ VPWR VGND sg13g2_nor2_1
XFILLER_22_988 VPWR VGND sg13g2_decap_8
X_4758_ net686 net734 _0188_ VPWR VGND sg13g2_nor2_1
X_3709_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[2\] net556 _1378_ VPWR
+ VGND sg13g2_nor2_1
X_4689_ net675 net727 _0119_ VPWR VGND sg13g2_nor2_1
XFILLER_1_837 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_0_358 VPWR VGND sg13g2_decap_4
XFILLER_1_1019 VPWR VGND sg13g2_decap_8
XFILLER_17_74 VPWR VGND sg13g2_fill_1
XFILLER_13_933 VPWR VGND sg13g2_decap_8
XFILLER_33_51 VPWR VGND sg13g2_fill_2
XFILLER_40_785 VPWR VGND sg13g2_decap_8
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_8_447 VPWR VGND sg13g2_decap_4
XFILLER_12_498 VPWR VGND sg13g2_decap_8
X_5175__74 VPWR VGND net74 sg13g2_tiehi
Xhold3 serialize.n420\[2\] VPWR VGND net408 sg13g2_dlygate4sd3_1
XFILLER_48_830 VPWR VGND sg13g2_decap_8
XFILLER_35_502 VPWR VGND sg13g2_decap_4
X_3991_ _1658_ VPWR _1659_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[0\]
+ net554 sg13g2_o21ai_1
XFILLER_22_229 VPWR VGND sg13g2_decap_4
X_2942_ VGND VPWR _0635_ _0786_ _0398_ _0788_ sg13g2_a21oi_1
XFILLER_30_240 VPWR VGND sg13g2_decap_8
X_2873_ _0685_ VPWR _0770_ VGND _0693_ _0695_ sg13g2_o21ai_1
XFILLER_30_251 VPWR VGND sg13g2_fill_2
X_4612_ net689 net739 _0042_ VPWR VGND sg13g2_nor2_1
X_4543_ tmds_blue.n193 _2136_ net603 _2172_ VPWR VGND sg13g2_nand3_1
X_4474_ _2090_ _2107_ _2080_ _2108_ VPWR VGND sg13g2_nand3_1
X_3425_ _1067_ _1068_ _1093_ _1094_ VPWR VGND sg13g2_nor3_1
X_3356_ _1038_ net797 _1037_ VPWR VGND sg13g2_nand2_1
X_3287_ _0643_ _0942_ _0981_ VPWR VGND sg13g2_nor2_2
X_5026_ net192 VGND VPWR _0454_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[1\]
+ _0111_ sg13g2_dfrbpq_1
XFILLER_21_240 VPWR VGND sg13g2_fill_1
XFILLER_21_251 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_10_958 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_decap_8
XFILLER_49_649 VPWR VGND sg13g2_fill_2
XFILLER_49_627 VPWR VGND sg13g2_decap_4
XFILLER_48_159 VPWR VGND sg13g2_fill_2
XFILLER_17_535 VPWR VGND sg13g2_decap_8
XFILLER_17_579 VPWR VGND sg13g2_decap_8
XFILLER_12_262 VPWR VGND sg13g2_fill_1
XFILLER_9_767 VPWR VGND sg13g2_fill_2
XFILLER_8_299 VPWR VGND sg13g2_decap_8
XFILLER_5_951 VPWR VGND sg13g2_decap_8
XFILLER_5_55 VPWR VGND sg13g2_fill_1
XFILLER_5_44 VPWR VGND sg13g2_decap_8
XFILLER_4_461 VPWR VGND sg13g2_fill_1
X_3210_ videogen.fancy_shader.video_x\[6\] _0815_ _0929_ VPWR VGND sg13g2_nor2_1
X_4190_ _1852_ _1840_ _1845_ VPWR VGND sg13g2_nand2_1
X_3141_ VGND VPWR tmds_red.n126 tmds_red.n132 _0870_ tmds_red.n100 sg13g2_a21oi_1
X_5081__371 VPWR VGND net371 sg13g2_tiehi
X_3072_ serialize.n452 serialize.n450 clknet_1_1__leaf_clk net6 VPWR VGND sg13g2_mux2_1
XFILLER_36_800 VPWR VGND sg13g2_fill_1
XFILLER_35_343 VPWR VGND sg13g2_fill_2
XFILLER_23_538 VPWR VGND sg13g2_fill_2
X_3974_ net612 _1630_ _1641_ _1642_ VPWR VGND sg13g2_nor3_2
X_2925_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\] _0783_ _0410_
+ VPWR VGND sg13g2_mux2_1
X_2856_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[0\] net790 _0764_ _0461_
+ VPWR VGND sg13g2_mux2_1
X_2787_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\] net774 _0749_ _0523_
+ VPWR VGND sg13g2_mux2_1
X_4526_ net602 _2152_ _2156_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
X_4457_ _2090_ _2091_ _2092_ VPWR VGND sg13g2_nor2_1
Xfanout702 net703 net702 VPWR VGND sg13g2_buf_8
X_3408_ _1074_ _1075_ _1077_ VPWR VGND sg13g2_and2_1
Xfanout724 net744 net724 VPWR VGND sg13g2_buf_8
Xfanout713 net714 net713 VPWR VGND sg13g2_buf_1
Xfanout735 net738 net735 VPWR VGND sg13g2_buf_1
Xfanout746 net751 net746 VPWR VGND sg13g2_buf_8
Xfanout757 net761 net757 VPWR VGND sg13g2_buf_8
X_4388_ _2032_ _2024_ _2033_ VPWR VGND sg13g2_xor2_1
X_5008__228 VPWR VGND net228 sg13g2_tiehi
X_3339_ _0642_ _1023_ _1026_ VPWR VGND sg13g2_nor2_1
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
Xfanout779 net783 net779 VPWR VGND sg13g2_buf_8
X_5009_ net226 VGND VPWR _0437_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[0\]
+ _0094_ sg13g2_dfrbpq_1
XFILLER_41_324 VPWR VGND sg13g2_fill_1
XFILLER_41_302 VPWR VGND sg13g2_decap_4
XFILLER_14_42 VPWR VGND sg13g2_decap_8
XFILLER_10_722 VPWR VGND sg13g2_fill_1
XFILLER_14_86 VPWR VGND sg13g2_fill_1
XFILLER_6_737 VPWR VGND sg13g2_decap_4
XFILLER_5_236 VPWR VGND sg13g2_fill_1
XFILLER_2_943 VPWR VGND sg13g2_decap_8
X_5130__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_17_310 VPWR VGND sg13g2_fill_1
XFILLER_45_663 VPWR VGND sg13g2_decap_8
XFILLER_17_376 VPWR VGND sg13g2_fill_2
XFILLER_17_398 VPWR VGND sg13g2_fill_2
XFILLER_20_508 VPWR VGND sg13g2_fill_1
XFILLER_20_519 VPWR VGND sg13g2_decap_8
X_2710_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[2\] net770 _0729_ _0580_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_553 VPWR VGND sg13g2_fill_1
X_3690_ _1355_ _1356_ _1357_ _1358_ _1359_ VPWR VGND sg13g2_nor4_1
X_4855__129 VPWR VGND net129 sg13g2_tiehi
X_2641_ _0694_ _0692_ VPWR VGND net610 sg13g2_nand2b_2
X_4311_ _1973_ _0662_ _1591_ VPWR VGND sg13g2_nand2_1
X_4242_ _1894_ _1900_ _1902_ _1904_ VPWR VGND sg13g2_or3_1
X_4173_ _1820_ _1827_ _1830_ _1835_ VPWR VGND sg13g2_or3_1
XFILLER_49_980 VPWR VGND sg13g2_decap_8
X_3124_ _0654_ net571 _0271_ VPWR VGND sg13g2_nor2_1
X_3055_ _0841_ _0648_ _0837_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_118 VPWR VGND sg13g2_fill_1
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
X_3957_ net618 VPWR _1625_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\]
+ net550 sg13g2_o21ai_1
X_2908_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[2\] net765 _0779_ _0423_
+ VPWR VGND sg13g2_mux2_1
Xclkbuf_0_clk_regs clk_regs clknet_0_clk_regs VPWR VGND sg13g2_buf_8
X_3888_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\] net550 _1557_ VPWR
+ VGND sg13g2_nor2_1
X_2839_ net780 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[1\] _0761_ _0474_
+ VPWR VGND sg13g2_mux2_1
X_4509_ tmds_blue.n193 tmds_blue.n132 _2139_ VPWR VGND sg13g2_xor2_1
XFILLER_4_8 VPWR VGND sg13g2_decap_8
XFILLER_47_906 VPWR VGND sg13g2_decap_8
Xfanout554 net555 net554 VPWR VGND sg13g2_buf_8
Xfanout565 _1303_ net565 VPWR VGND sg13g2_buf_8
XFILLER_19_619 VPWR VGND sg13g2_fill_1
Xfanout587 _0687_ net587 VPWR VGND sg13g2_buf_8
Xfanout598 _0645_ net598 VPWR VGND sg13g2_buf_8
Xfanout576 net577 net576 VPWR VGND sg13g2_buf_8
XFILLER_27_630 VPWR VGND sg13g2_fill_2
XFILLER_42_655 VPWR VGND sg13g2_fill_2
XFILLER_26_195 VPWR VGND sg13g2_decap_8
XFILLER_10_574 VPWR VGND sg13g2_decap_8
XFILLER_49_265 VPWR VGND sg13g2_decap_4
XFILLER_46_972 VPWR VGND sg13g2_decap_8
XFILLER_18_696 VPWR VGND sg13g2_fill_1
X_4860_ net119 VGND VPWR _0288_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\]
+ _0019_ sg13g2_dfrbpq_1
X_3811_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\] net557 _1480_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_143 VPWR VGND sg13g2_fill_1
X_4791_ net690 net742 _0221_ VPWR VGND sg13g2_nor2_1
X_3742_ net622 VPWR _1411_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[1\]
+ net555 sg13g2_o21ai_1
XFILLER_9_383 VPWR VGND sg13g2_fill_2
X_3673_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[2\] net586 _1342_ VPWR
+ VGND sg13g2_nor2_1
X_2624_ _0675_ _0676_ _0677_ VPWR VGND sg13g2_and2_1
X_4225_ _1887_ _1803_ _1878_ VPWR VGND sg13g2_xnor2_1
X_4156_ VPWR VGND _1811_ _1805_ _1817_ _1812_ _1818_ _1813_ sg13g2_a221oi_1
X_3107_ net426 red_tmds_par\[5\] net696 serialize.n427\[5\] VPWR VGND sg13g2_mux2_1
X_4087_ _1741_ _1751_ _1752_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_972 VPWR VGND sg13g2_decap_8
X_3038_ VGND VPWR net595 net11 _0690_ net549 sg13g2_a21oi_2
XFILLER_24_633 VPWR VGND sg13g2_decap_8
XFILLER_24_644 VPWR VGND sg13g2_fill_2
XFILLER_36_493 VPWR VGND sg13g2_fill_1
XFILLER_23_154 VPWR VGND sg13g2_fill_2
X_4989_ net269 VGND VPWR _0417_ videogen.test_lut_thingy.pixel_feeder_inst.row\[55\]\[0\]
+ _0074_ sg13g2_dfrbpq_1
XFILLER_23_176 VPWR VGND sg13g2_decap_8
XFILLER_3_515 VPWR VGND sg13g2_fill_1
XFILLER_19_416 VPWR VGND sg13g2_decap_4
XFILLER_28_950 VPWR VGND sg13g2_decap_8
XFILLER_36_73 VPWR VGND sg13g2_fill_1
XFILLER_43_997 VPWR VGND sg13g2_decap_8
XFILLER_14_154 VPWR VGND sg13g2_decap_4
XFILLER_15_655 VPWR VGND sg13g2_decap_8
X_5136__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_7_810 VPWR VGND sg13g2_fill_1
XFILLER_6_375 VPWR VGND sg13g2_fill_2
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
X_4010_ net596 _1672_ _1677_ _1678_ VPWR VGND sg13g2_nor3_1
XFILLER_26_909 VPWR VGND sg13g2_decap_8
XFILLER_18_460 VPWR VGND sg13g2_fill_1
XFILLER_19_972 VPWR VGND sg13g2_decap_8
X_4912_ net398 VGND VPWR _0340_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[2\]
+ _0040_ sg13g2_dfrbpq_1
XFILLER_34_964 VPWR VGND sg13g2_decap_8
X_4843_ net145 VGND VPWR _0271_ green_tmds_par\[0\] net643 sg13g2_dfrbpq_1
XFILLER_21_647 VPWR VGND sg13g2_fill_1
X_4774_ net658 net710 _0204_ VPWR VGND sg13g2_nor2_1
XFILLER_21_658 VPWR VGND sg13g2_decap_8
X_3725_ net611 _1382_ _1393_ _1394_ VPWR VGND sg13g2_nor3_1
X_5154__297 VPWR VGND net297 sg13g2_tiehi
X_3656_ net598 VPWR _1325_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\]
+ net551 sg13g2_o21ai_1
X_3587_ _1166_ VPWR _1256_ VGND _1138_ _1158_ sg13g2_o21ai_1
X_2607_ VPWR _0663_ tmds_red.n102 VGND sg13g2_inv_1
XFILLER_0_529 VPWR VGND sg13g2_decap_8
X_4208_ _1870_ _1192_ _1869_ VPWR VGND sg13g2_nand2_2
X_5188_ net211 VGND VPWR _0612_ blue_tmds_par\[2\] net637 sg13g2_dfrbpq_1
X_4139_ _1757_ _1011_ _1801_ VPWR VGND sg13g2_xor2_1
XFILLER_43_205 VPWR VGND sg13g2_fill_2
XFILLER_43_249 VPWR VGND sg13g2_decap_8
XFILLER_25_942 VPWR VGND sg13g2_decap_8
XFILLER_40_901 VPWR VGND sg13g2_decap_4
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_7_128 VPWR VGND sg13g2_decap_8
XFILLER_11_157 VPWR VGND sg13g2_fill_1
XFILLER_4_813 VPWR VGND sg13g2_decap_8
XFILLER_26_1007 VPWR VGND sg13g2_decap_8
XFILLER_16_931 VPWR VGND sg13g2_decap_8
XFILLER_30_422 VPWR VGND sg13g2_fill_2
XFILLER_31_956 VPWR VGND sg13g2_decap_8
X_3510_ _1077_ _1170_ _1178_ _1179_ VPWR VGND sg13g2_nor3_1
X_4490_ _2123_ _2077_ _2090_ VPWR VGND sg13g2_nand2_1
X_3441_ _1107_ _1109_ _1092_ _1110_ VPWR VGND sg13g2_nand3_1
X_3372_ _0673_ _1043_ _1049_ VPWR VGND sg13g2_nor2_1
X_5149__377 VPWR VGND net377 sg13g2_tiehi
X_5111_ net244 VGND VPWR _0535_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[1\]
+ _0183_ sg13g2_dfrbpq_1
X_5042_ net160 VGND VPWR _0470_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[1\]
+ _0127_ sg13g2_dfrbpq_1
XFILLER_26_717 VPWR VGND sg13g2_decap_4
XFILLER_41_709 VPWR VGND sg13g2_decap_8
XFILLER_34_761 VPWR VGND sg13g2_fill_1
X_4921__380 VPWR VGND net380 sg13g2_tiehi
X_4826_ net657 net709 _0256_ VPWR VGND sg13g2_nor2_1
XFILLER_22_967 VPWR VGND sg13g2_decap_8
X_4757_ net683 net734 _0187_ VPWR VGND sg13g2_nor2_1
X_3708_ net616 VPWR _1377_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\]
+ net588 sg13g2_o21ai_1
X_4688_ net676 net728 _0118_ VPWR VGND sg13g2_nor2_1
X_3639_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\] net581 _1308_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_1_816 VPWR VGND sg13g2_decap_8
X_5204__316 VPWR VGND net316 sg13g2_tiehi
X_5126__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_44_558 VPWR VGND sg13g2_fill_2
XFILLER_17_86 VPWR VGND sg13g2_decap_8
XFILLER_13_912 VPWR VGND sg13g2_decap_8
XFILLER_12_422 VPWR VGND sg13g2_decap_8
XFILLER_33_41 VPWR VGND sg13g2_fill_1
X_5018__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_13_989 VPWR VGND sg13g2_decap_8
XFILLER_4_621 VPWR VGND sg13g2_decap_8
Xhold4 serialize.n420\[3\] VPWR VGND net409 sg13g2_dlygate4sd3_1
XFILLER_48_886 VPWR VGND sg13g2_decap_8
X_3990_ _1658_ net594 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
X_2941_ net776 _0786_ _0788_ VPWR VGND sg13g2_nor2_1
X_4611_ net655 net707 _0041_ VPWR VGND sg13g2_nor2_1
X_2872_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\] _0768_ _0449_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_982 VPWR VGND sg13g2_decap_8
X_4542_ VGND VPWR _2164_ _2168_ _2171_ _2170_ sg13g2_a21oi_1
X_4473_ _2107_ _2104_ _2105_ VPWR VGND sg13g2_xnor2_1
X_3424_ VGND VPWR _1093_ _1085_ _1070_ sg13g2_or2_1
X_3355_ _1035_ _1036_ _0922_ _1037_ VPWR VGND sg13g2_nand3_1
X_3286_ _0975_ _0980_ _0337_ VPWR VGND sg13g2_nor2_1
X_4865__109 VPWR VGND net109 sg13g2_tiehi
X_5025_ net194 VGND VPWR _0453_ videogen.test_lut_thingy.pixel_feeder_inst.row\[46\]\[0\]
+ _0110_ sg13g2_dfrbpq_1
XFILLER_38_341 VPWR VGND sg13g2_fill_2
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
XFILLER_10_937 VPWR VGND sg13g2_decap_8
XFILLER_22_786 VPWR VGND sg13g2_decap_8
X_5052__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_22_797 VPWR VGND sg13g2_fill_2
X_4809_ net689 net739 _0239_ VPWR VGND sg13g2_nor2_1
X_4904__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_0_101 VPWR VGND sg13g2_decap_4
XFILLER_28_41 VPWR VGND sg13g2_decap_8
XFILLER_45_867 VPWR VGND sg13g2_fill_1
XFILLER_44_399 VPWR VGND sg13g2_fill_2
XFILLER_8_212 VPWR VGND sg13g2_fill_1
XFILLER_8_223 VPWR VGND sg13g2_fill_2
XFILLER_9_746 VPWR VGND sg13g2_fill_1
XFILLER_8_278 VPWR VGND sg13g2_decap_8
XFILLER_5_930 VPWR VGND sg13g2_decap_8
X_3140_ _0869_ tmds_red.n114 tmds_red.n132 VPWR VGND sg13g2_xnor2_1
X_3071_ serialize.n455 serialize.n453 clknet_1_1__leaf_clk net5 VPWR VGND sg13g2_mux2_1
XFILLER_36_823 VPWR VGND sg13g2_fill_1
XFILLER_36_878 VPWR VGND sg13g2_decap_8
X_3973_ net614 _1635_ _1640_ _1641_ VPWR VGND sg13g2_nor3_1
X_2924_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\] _0783_ _0411_
+ VPWR VGND sg13g2_mux2_1
X_2855_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[1\] net779 _0764_ _0462_
+ VPWR VGND sg13g2_mux2_1
X_4525_ _2155_ net602 _2154_ VPWR VGND sg13g2_nand2_1
X_2786_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\] net767 _0749_ _0524_
+ VPWR VGND sg13g2_mux2_1
X_5139__86 VPWR VGND net86 sg13g2_tiehi
X_4456_ _0857_ VPWR _2091_ VGND tmds_green.dc_balancing_reg\[1\] _0858_ sg13g2_o21ai_1
Xfanout703 net706 net703 VPWR VGND sg13g2_buf_8
X_3407_ _1076_ _1074_ _1075_ VPWR VGND sg13g2_nand2_2
Xfanout714 net724 net714 VPWR VGND sg13g2_buf_8
X_4387_ _1998_ VPWR _2032_ VGND _0903_ _0905_ sg13g2_o21ai_1
Xfanout736 net737 net736 VPWR VGND sg13g2_buf_8
X_3338_ _0642_ _1023_ _1025_ VPWR VGND sg13g2_and2_1
Xfanout725 net726 net725 VPWR VGND sg13g2_buf_8
Xfanout758 net761 net758 VPWR VGND sg13g2_buf_8
Xfanout747 net748 net747 VPWR VGND sg13g2_buf_8
Xfanout769 net772 net769 VPWR VGND sg13g2_buf_8
X_3269_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[1\] _0968_ _0970_ VPWR
+ VGND sg13g2_nor2_1
X_5008_ net228 VGND VPWR _0436_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[3\]
+ _0093_ sg13g2_dfrbpq_1
XFILLER_27_867 VPWR VGND sg13g2_decap_4
XFILLER_10_767 VPWR VGND sg13g2_fill_2
XFILLER_30_20 VPWR VGND sg13g2_fill_2
XFILLER_2_922 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_999 VPWR VGND sg13g2_decap_8
XFILLER_49_458 VPWR VGND sg13g2_decap_8
XFILLER_49_425 VPWR VGND sg13g2_decap_8
XFILLER_39_62 VPWR VGND sg13g2_fill_1
XFILLER_45_631 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
X_2640_ _0693_ net611 _0689_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_771 VPWR VGND sg13g2_decap_8
X_4310_ _1972_ _1963_ _1971_ VPWR VGND sg13g2_nand2_1
X_4241_ _1903_ _1899_ _1902_ VPWR VGND sg13g2_nand2b_1
X_4172_ VGND VPWR _1834_ _1830_ _1827_ sg13g2_or2_1
X_3123_ _0266_ net796 net739 net432 VPWR VGND sg13g2_and3_1
X_3054_ _0648_ _0837_ _0840_ VPWR VGND sg13g2_nor2_2
XFILLER_36_620 VPWR VGND sg13g2_fill_1
X_3956_ net618 _1620_ _1621_ _1623_ _1624_ VPWR VGND sg13g2_nor4_1
XFILLER_11_509 VPWR VGND sg13g2_decap_8
X_2907_ videogen.test_lut_thingy.pixel_feeder_inst.row\[54\]\[3\] net755 _0779_ _0424_
+ VPWR VGND sg13g2_mux2_1
X_5157__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_32_881 VPWR VGND sg13g2_fill_2
X_3887_ videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\] net573 _1556_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_31_391 VPWR VGND sg13g2_decap_4
X_2838_ net768 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[2\] _0761_ _0475_
+ VPWR VGND sg13g2_mux2_1
X_2769_ _0746_ _0720_ _0744_ VPWR VGND sg13g2_nand2_2
X_4508_ VGND VPWR _2065_ _2136_ _2138_ _2137_ sg13g2_a21oi_1
X_4439_ _2076_ net801 _2075_ VPWR VGND sg13g2_nand2_1
Xfanout544 _1089_ net544 VPWR VGND sg13g2_buf_8
Xfanout566 net567 net566 VPWR VGND sg13g2_buf_8
Xfanout555 _1300_ net555 VPWR VGND sg13g2_buf_8
X_4886__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_46_406 VPWR VGND sg13g2_decap_8
Xfanout599 tmds_green.n132 net599 VPWR VGND sg13g2_buf_8
Xfanout577 _0702_ net577 VPWR VGND sg13g2_buf_8
Xfanout588 net592 net588 VPWR VGND sg13g2_buf_8
XFILLER_18_119 VPWR VGND sg13g2_decap_4
X_5205__285 VPWR VGND net285 sg13g2_tiehi
XFILLER_15_804 VPWR VGND sg13g2_fill_1
XFILLER_41_111 VPWR VGND sg13g2_fill_1
XFILLER_25_42 VPWR VGND sg13g2_decap_8
X_5063__55 VPWR VGND net55 sg13g2_tiehi
XFILLER_25_86 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_10_531 VPWR VGND sg13g2_fill_2
XFILLER_6_524 VPWR VGND sg13g2_fill_2
XFILLER_2_796 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_46_951 VPWR VGND sg13g2_decap_8
XFILLER_17_174 VPWR VGND sg13g2_decap_8
XFILLER_17_196 VPWR VGND sg13g2_decap_8
XFILLER_32_100 VPWR VGND sg13g2_decap_4
XFILLER_33_656 VPWR VGND sg13g2_decap_4
X_4790_ net685 net737 _0220_ VPWR VGND sg13g2_nor2_1
X_3810_ net596 _1473_ _1478_ _1479_ VPWR VGND sg13g2_nor3_1
XFILLER_20_306 VPWR VGND sg13g2_fill_1
XFILLER_33_678 VPWR VGND sg13g2_decap_8
X_3741_ net617 _1404_ _1409_ _1410_ VPWR VGND sg13g2_nor3_1
X_3672_ net598 VPWR _1341_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\]
+ net562 sg13g2_o21ai_1
X_2623_ videogen.fancy_shader.video_y\[3\] videogen.fancy_shader.video_y\[2\] videogen.fancy_shader.video_y\[1\]
+ net608 _0676_ VPWR VGND sg13g2_nor4_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_4224_ _1886_ _1147_ _1885_ VPWR VGND sg13g2_xnor2_1
X_4155_ _1808_ _1811_ _1804_ _1817_ VPWR VGND _1813_ sg13g2_nand4_1
X_3106_ net442 red_tmds_par\[4\] net696 serialize.n427\[4\] VPWR VGND sg13g2_mux2_1
X_4086_ _1738_ VPWR _1751_ VGND _1734_ _1740_ sg13g2_o21ai_1
X_3037_ VGND VPWR net595 net10 _0709_ net549 sg13g2_a21oi_2
XFILLER_24_612 VPWR VGND sg13g2_decap_8
X_4988_ net270 VGND VPWR _0416_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\]
+ _0073_ sg13g2_dfrbpq_1
XFILLER_11_306 VPWR VGND sg13g2_decap_8
X_3939_ net617 _1601_ _1606_ _1607_ VPWR VGND sg13g2_nor3_1
X_4931__360 VPWR VGND net360 sg13g2_tiehi
XFILLER_46_214 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_fill_1
XFILLER_36_30 VPWR VGND sg13g2_fill_2
XFILLER_14_111 VPWR VGND sg13g2_fill_1
XFILLER_43_976 VPWR VGND sg13g2_decap_8
XFILLER_42_464 VPWR VGND sg13g2_decap_4
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_14_199 VPWR VGND sg13g2_fill_2
XFILLER_11_862 VPWR VGND sg13g2_fill_2
XFILLER_7_899 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_4
XFILLER_2_560 VPWR VGND sg13g2_decap_8
XFILLER_38_704 VPWR VGND sg13g2_fill_1
XFILLER_28_5 VPWR VGND sg13g2_fill_2
X_5108__256 VPWR VGND net256 sg13g2_tiehi
XFILLER_19_951 VPWR VGND sg13g2_decap_8
X_4911_ net400 VGND VPWR _0339_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[1\]
+ _0039_ sg13g2_dfrbpq_1
XFILLER_18_472 VPWR VGND sg13g2_fill_2
XFILLER_34_943 VPWR VGND sg13g2_decap_8
X_4842_ net147 VGND VPWR _0270_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[3\]
+ _0009_ sg13g2_dfrbpq_1
X_4773_ net667 net720 _0203_ VPWR VGND sg13g2_nor2_1
X_3724_ net623 _1387_ _1392_ _1393_ VPWR VGND sg13g2_nor3_1
X_3655_ net613 VPWR _1324_ VGND _1317_ _1323_ sg13g2_o21ai_1
X_2606_ _0662_ net1 VPWR VGND sg13g2_inv_2
X_3586_ _1255_ _1248_ _1251_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_508 VPWR VGND sg13g2_decap_8
X_4207_ _0994_ _1059_ _1869_ VPWR VGND sg13g2_nor2b_2
XFILLER_29_704 VPWR VGND sg13g2_fill_2
X_5187_ net219 VGND VPWR _0611_ blue_tmds_par\[1\] net643 sg13g2_dfrbpq_1
XFILLER_29_715 VPWR VGND sg13g2_fill_1
X_4138_ _1012_ _1011_ _1800_ VPWR VGND sg13g2_xor2_1
XFILLER_44_729 VPWR VGND sg13g2_fill_2
X_4069_ _1733_ VPWR _1734_ VGND _1726_ _1730_ sg13g2_o21ai_1
XFILLER_25_921 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_24_497 VPWR VGND sg13g2_decap_4
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_8_608 VPWR VGND sg13g2_fill_2
XFILLER_20_670 VPWR VGND sg13g2_decap_8
XFILLER_3_302 VPWR VGND sg13g2_decap_8
XFILLER_22_98 VPWR VGND sg13g2_decap_8
XFILLER_4_869 VPWR VGND sg13g2_decap_8
XFILLER_3_346 VPWR VGND sg13g2_fill_1
XFILLER_47_51 VPWR VGND sg13g2_decap_8
XFILLER_47_589 VPWR VGND sg13g2_decap_8
XFILLER_16_910 VPWR VGND sg13g2_decap_8
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_43_773 VPWR VGND sg13g2_fill_2
XFILLER_31_935 VPWR VGND sg13g2_decap_8
XFILLER_11_692 VPWR VGND sg13g2_fill_2
XFILLER_6_184 VPWR VGND sg13g2_decap_8
X_3440_ videogen.fancy_shader.n646\[9\] videogen.fancy_shader.video_y\[9\] _1109_
+ VPWR VGND sg13g2_xor2_1
X_3371_ VGND VPWR videogen.fancy_shader.video_y\[6\] _1046_ _1048_ videogen.fancy_shader.video_y\[7\]
+ sg13g2_a21oi_1
X_5110_ net248 VGND VPWR _0534_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[0\]
+ _0182_ sg13g2_dfrbpq_1
X_5184__258 VPWR VGND net258 sg13g2_tiehi
X_5041_ net162 VGND VPWR _0469_ videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[0\]
+ _0126_ sg13g2_dfrbpq_1
XFILLER_19_792 VPWR VGND sg13g2_decap_8
XFILLER_34_740 VPWR VGND sg13g2_decap_8
XFILLER_34_751 VPWR VGND sg13g2_fill_1
X_4825_ net656 net708 _0255_ VPWR VGND sg13g2_nor2_1
XFILLER_22_946 VPWR VGND sg13g2_decap_8
XFILLER_21_489 VPWR VGND sg13g2_fill_1
X_4756_ net683 net735 _0186_ VPWR VGND sg13g2_nor2_1
X_3707_ _1372_ _1373_ _1374_ _1375_ _1376_ VPWR VGND sg13g2_nor4_1
X_4687_ net676 net728 _0117_ VPWR VGND sg13g2_nor2_1
XFILLER_49_1008 VPWR VGND sg13g2_decap_8
X_3638_ net597 VPWR _1307_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\]
+ net559 sg13g2_o21ai_1
X_3569_ VGND VPWR _1222_ _1229_ _1238_ _1237_ sg13g2_a21oi_1
XFILLER_0_338 VPWR VGND sg13g2_fill_1
XFILLER_0_349 VPWR VGND sg13g2_decap_4
X_5239_ net805 VGND VPWR serialize.n427\[0\] serialize.n450 clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_17_718 VPWR VGND sg13g2_decap_8
XFILLER_12_401 VPWR VGND sg13g2_decap_8
XFILLER_25_773 VPWR VGND sg13g2_decap_4
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_13_968 VPWR VGND sg13g2_decap_8
XFILLER_24_283 VPWR VGND sg13g2_fill_1
XFILLER_33_31 VPWR VGND sg13g2_fill_1
XFILLER_12_478 VPWR VGND sg13g2_decap_8
XFILLER_33_97 VPWR VGND sg13g2_decap_8
XFILLER_39_309 VPWR VGND sg13g2_decap_8
Xhold5 serialize.n420\[0\] VPWR VGND net410 sg13g2_dlygate4sd3_1
XFILLER_47_331 VPWR VGND sg13g2_decap_4
XFILLER_0_894 VPWR VGND sg13g2_decap_8
XFILLER_48_865 VPWR VGND sg13g2_decap_8
XFILLER_35_515 VPWR VGND sg13g2_decap_8
XFILLER_16_762 VPWR VGND sg13g2_decap_4
X_2940_ VGND VPWR _0634_ _0786_ _0399_ _0787_ sg13g2_a21oi_1
X_2871_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\] _0768_ _0450_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_732 VPWR VGND sg13g2_decap_8
X_4610_ net655 net707 _0040_ VPWR VGND sg13g2_nor2_1
XFILLER_8_961 VPWR VGND sg13g2_decap_8
X_4541_ VGND VPWR _2151_ _2153_ _2170_ _2169_ sg13g2_a21oi_1
X_4472_ _2106_ _2104_ _2105_ VPWR VGND sg13g2_nand2b_1
XFILLER_7_471 VPWR VGND sg13g2_fill_2
X_3423_ _1092_ videogen.fancy_shader.video_y\[8\] net609 VPWR VGND sg13g2_nand2_1
X_3354_ _0637_ videogen.fancy_shader.video_y\[8\] _0831_ _0935_ _1036_ VPWR VGND sg13g2_nor4_1
XFILLER_31_0 VPWR VGND sg13g2_decap_8
X_3285_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] _0977_
+ _0980_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] sg13g2_a21oi_1
XFILLER_38_331 VPWR VGND sg13g2_decap_4
X_5024_ net196 VGND VPWR _0452_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[3\]
+ _0109_ sg13g2_dfrbpq_1
XFILLER_10_916 VPWR VGND sg13g2_decap_8
X_4808_ net688 net740 _0238_ VPWR VGND sg13g2_nor2_1
X_4739_ net678 net732 _0169_ VPWR VGND sg13g2_nor2_1
XFILLER_0_135 VPWR VGND sg13g2_decap_4
XFILLER_0_179 VPWR VGND sg13g2_decap_4
XFILLER_28_20 VPWR VGND sg13g2_decap_8
XFILLER_28_75 VPWR VGND sg13g2_decap_4
XFILLER_44_312 VPWR VGND sg13g2_decap_8
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_25_570 VPWR VGND sg13g2_fill_2
XFILLER_32_507 VPWR VGND sg13g2_fill_1
XFILLER_32_529 VPWR VGND sg13g2_fill_1
XFILLER_44_63 VPWR VGND sg13g2_fill_1
XFILLER_13_721 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_40_595 VPWR VGND sg13g2_decap_8
XFILLER_9_769 VPWR VGND sg13g2_fill_1
XFILLER_12_275 VPWR VGND sg13g2_decap_8
XFILLER_8_257 VPWR VGND sg13g2_fill_2
XFILLER_4_452 VPWR VGND sg13g2_decap_8
XFILLER_5_986 VPWR VGND sg13g2_decap_8
XFILLER_4_496 VPWR VGND sg13g2_decap_8
X_3070_ serialize.n458 serialize.n456 clknet_1_0__leaf_clk net3 VPWR VGND sg13g2_mux2_1
XFILLER_0_691 VPWR VGND sg13g2_decap_8
XFILLER_39_1018 VPWR VGND sg13g2_decap_8
XFILLER_35_345 VPWR VGND sg13g2_fill_1
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_3972_ net621 _1636_ _1637_ _1639_ _1640_ VPWR VGND sg13g2_nor4_1
X_2923_ net755 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\] _0783_ _0412_
+ VPWR VGND sg13g2_mux2_1
X_2854_ videogen.test_lut_thingy.pixel_feeder_inst.row\[44\]\[2\] net767 _0764_ _0463_
+ VPWR VGND sg13g2_mux2_1
X_2785_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\] net752 _0749_ _0525_
+ VPWR VGND sg13g2_mux2_1
X_4524_ _2152_ _2134_ _2154_ VPWR VGND sg13g2_xor2_1
X_4455_ _2090_ tmds_green.dc_balancing_reg\[2\] _2088_ VPWR VGND sg13g2_xnor2_1
Xfanout715 net718 net715 VPWR VGND sg13g2_buf_8
X_3406_ _1075_ _1009_ _1073_ VPWR VGND sg13g2_nand2_1
Xfanout704 net705 net704 VPWR VGND sg13g2_buf_8
X_4386_ VGND VPWR _2000_ _2011_ _2031_ _2013_ sg13g2_a21oi_1
Xfanout737 net738 net737 VPWR VGND sg13g2_buf_8
X_3337_ _1022_ _1024_ _0352_ VPWR VGND sg13g2_nor2_1
Xfanout726 net733 net726 VPWR VGND sg13g2_buf_8
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_8
Xfanout759 net761 net759 VPWR VGND sg13g2_buf_8
XFILLER_39_640 VPWR VGND sg13g2_fill_1
X_3268_ _0967_ _0968_ _0969_ _0330_ VPWR VGND sg13g2_nor3_1
X_5007_ net230 VGND VPWR _0435_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[2\]
+ _0092_ sg13g2_dfrbpq_1
XFILLER_39_673 VPWR VGND sg13g2_fill_1
X_3199_ videogen.fancy_shader.video_x\[0\] _0923_ _0299_ VPWR VGND sg13g2_nor2_1
XFILLER_27_813 VPWR VGND sg13g2_fill_1
XFILLER_14_529 VPWR VGND sg13g2_decap_8
XFILLER_22_562 VPWR VGND sg13g2_decap_8
XFILLER_10_735 VPWR VGND sg13g2_fill_2
XFILLER_22_573 VPWR VGND sg13g2_fill_1
XFILLER_6_706 VPWR VGND sg13g2_decap_4
XFILLER_2_901 VPWR VGND sg13g2_decap_8
XFILLER_49_404 VPWR VGND sg13g2_decap_8
XFILLER_2_978 VPWR VGND sg13g2_decap_8
XFILLER_49_437 VPWR VGND sg13g2_decap_8
XFILLER_45_610 VPWR VGND sg13g2_fill_1
XFILLER_29_172 VPWR VGND sg13g2_decap_4
XFILLER_17_378 VPWR VGND sg13g2_fill_1
XFILLER_33_816 VPWR VGND sg13g2_decap_8
XFILLER_13_551 VPWR VGND sg13g2_decap_8
XFILLER_9_511 VPWR VGND sg13g2_fill_2
X_4240_ _1902_ _1828_ _1901_ VPWR VGND sg13g2_xnor2_1
X_4171_ _1823_ VPWR _1833_ VGND _1831_ _1832_ sg13g2_o21ai_1
X_3122_ VGND VPWR net739 net432 _0265_ _0854_ sg13g2_a21oi_1
X_5007__230 VPWR VGND net230 sg13g2_tiehi
X_3053_ VGND VPWR _0835_ _0839_ net14 _0836_ sg13g2_a21oi_1
XFILLER_27_109 VPWR VGND sg13g2_decap_8
XFILLER_23_304 VPWR VGND sg13g2_fill_2
XFILLER_35_186 VPWR VGND sg13g2_decap_8
X_3955_ _1622_ VPWR _1623_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[9\]\[0\]
+ net561 sg13g2_o21ai_1
X_2906_ _0707_ _0772_ _0779_ VPWR VGND sg13g2_nor2_2
X_3886_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[3\] net584 _1555_ VPWR
+ VGND sg13g2_nor2_1
X_2837_ net758 videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\] _0761_ _0476_
+ VPWR VGND sg13g2_mux2_1
X_2768_ _0745_ _0743_ VPWR VGND net545 sg13g2_nand2b_2
X_4918__386 VPWR VGND net386 sg13g2_tiehi
X_2699_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\] net775 _0725_ _0587_
+ VPWR VGND sg13g2_mux2_1
X_4507_ net603 _2071_ _2136_ _2137_ VPWR VGND sg13g2_nor3_1
X_4438_ _2075_ hsync tmds_blue.vsync VPWR VGND sg13g2_xnor2_1
X_5088__357 VPWR VGND net357 sg13g2_tiehi
Xfanout556 net560 net556 VPWR VGND sg13g2_buf_8
Xfanout545 _0691_ net545 VPWR VGND sg13g2_buf_8
X_4369_ net548 _0906_ _2015_ VPWR VGND sg13g2_nor2_1
Xfanout567 net570 net567 VPWR VGND sg13g2_buf_8
Xfanout589 net592 net589 VPWR VGND sg13g2_buf_8
Xfanout578 net582 net578 VPWR VGND sg13g2_buf_8
XFILLER_46_429 VPWR VGND sg13g2_decap_8
XFILLER_27_632 VPWR VGND sg13g2_fill_1
XFILLER_41_189 VPWR VGND sg13g2_decap_8
X_4854__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_775 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_4
XFILLER_49_234 VPWR VGND sg13g2_decap_8
XFILLER_18_610 VPWR VGND sg13g2_decap_4
XFILLER_46_930 VPWR VGND sg13g2_decap_8
XFILLER_17_120 VPWR VGND sg13g2_decap_4
XFILLER_17_153 VPWR VGND sg13g2_fill_2
XFILLER_33_613 VPWR VGND sg13g2_decap_8
XFILLER_33_635 VPWR VGND sg13g2_decap_8
X_3740_ net626 _1405_ _1406_ _1408_ _1409_ VPWR VGND sg13g2_nor4_1
XFILLER_13_381 VPWR VGND sg13g2_fill_1
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_3671_ _1336_ _1337_ _1338_ _1339_ _1340_ VPWR VGND sg13g2_nor4_1
X_2622_ videogen.fancy_shader.video_y\[4\] _0674_ _0675_ VPWR VGND sg13g2_nor2b_1
X_4223_ _1876_ _1802_ _1885_ VPWR VGND sg13g2_xor2_1
X_4154_ _1813_ VPWR _1816_ VGND _1807_ _1811_ sg13g2_o21ai_1
X_3105_ net424 red_tmds_par\[3\] net696 serialize.n427\[3\] VPWR VGND sg13g2_mux2_1
X_4085_ _1750_ _1748_ _1749_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_429 VPWR VGND sg13g2_decap_8
X_3036_ VGND VPWR net549 _0703_ net9 net595 sg13g2_a21oi_1
XFILLER_23_156 VPWR VGND sg13g2_fill_1
XFILLER_24_679 VPWR VGND sg13g2_decap_4
X_4987_ net272 VGND VPWR _0415_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[2\]
+ _0072_ sg13g2_dfrbpq_1
XFILLER_20_852 VPWR VGND sg13g2_decap_8
X_3938_ net626 _1602_ _1603_ _1605_ _1606_ VPWR VGND sg13g2_nor4_1
X_3869_ _1534_ _1535_ _1536_ _1537_ _1538_ VPWR VGND sg13g2_nor4_1
XFILLER_11_67 VPWR VGND sg13g2_fill_2
X_5129__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_46_259 VPWR VGND sg13g2_decap_4
XFILLER_28_985 VPWR VGND sg13g2_decap_8
XFILLER_42_421 VPWR VGND sg13g2_decap_4
XFILLER_43_955 VPWR VGND sg13g2_decap_8
XFILLER_15_646 VPWR VGND sg13g2_decap_4
XFILLER_30_627 VPWR VGND sg13g2_decap_8
XFILLER_30_638 VPWR VGND sg13g2_fill_2
XFILLER_11_841 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_fill_2
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_10_373 VPWR VGND sg13g2_fill_2
XFILLER_11_896 VPWR VGND sg13g2_decap_8
XFILLER_7_878 VPWR VGND sg13g2_decap_8
XFILLER_6_388 VPWR VGND sg13g2_fill_2
XFILLER_37_215 VPWR VGND sg13g2_decap_4
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_46_771 VPWR VGND sg13g2_fill_1
X_4910_ net404 VGND VPWR _0338_ videogen.test_lut_thingy.pixel_feeder_inst.row\[12\]\[0\]
+ _0038_ sg13g2_dfrbpq_1
XFILLER_18_495 VPWR VGND sg13g2_fill_1
XFILLER_34_922 VPWR VGND sg13g2_decap_8
X_4841_ net149 VGND VPWR _0269_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\]
+ _0008_ sg13g2_dfrbpq_1
XFILLER_33_443 VPWR VGND sg13g2_decap_8
XFILLER_21_638 VPWR VGND sg13g2_decap_8
XFILLER_33_476 VPWR VGND sg13g2_fill_1
XFILLER_34_999 VPWR VGND sg13g2_decap_8
X_4772_ net657 net709 _0202_ VPWR VGND sg13g2_nor2_1
X_3723_ _1388_ _1389_ _1390_ _1391_ _1392_ VPWR VGND sg13g2_nor4_1
XFILLER_9_182 VPWR VGND sg13g2_decap_8
X_3654_ net625 VPWR _1323_ VGND _1318_ _1322_ sg13g2_o21ai_1
X_2605_ _0661_ net2 VPWR VGND sg13g2_inv_2
X_3585_ _1247_ _1251_ _1146_ _1254_ VPWR VGND sg13g2_nand3_1
X_4206_ _1862_ VPWR _1868_ VGND _1866_ _1867_ sg13g2_o21ai_1
X_5186_ net227 VGND VPWR _0610_ blue_tmds_par\[0\] net637 sg13g2_dfrbpq_1
XFILLER_29_727 VPWR VGND sg13g2_decap_8
X_4137_ _1799_ _1694_ _1798_ VPWR VGND sg13g2_nand2b_1
X_4068_ _1726_ VPWR _1733_ VGND _1730_ _1731_ sg13g2_o21ai_1
XFILLER_25_900 VPWR VGND sg13g2_decap_8
XFILLER_37_782 VPWR VGND sg13g2_fill_1
X_3019_ videogen.fancy_shader.video_x\[5\] _0814_ _0815_ VPWR VGND sg13g2_and2_1
XFILLER_25_977 VPWR VGND sg13g2_decap_8
XFILLER_12_627 VPWR VGND sg13g2_fill_2
XFILLER_11_115 VPWR VGND sg13g2_decap_4
XFILLER_12_638 VPWR VGND sg13g2_decap_8
XFILLER_12_649 VPWR VGND sg13g2_decap_8
XFILLER_22_66 VPWR VGND sg13g2_decap_8
XFILLER_4_848 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_19_259 VPWR VGND sg13g2_decap_4
XFILLER_15_410 VPWR VGND sg13g2_fill_2
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_31_914 VPWR VGND sg13g2_decap_8
XFILLER_42_295 VPWR VGND sg13g2_fill_1
XFILLER_42_284 VPWR VGND sg13g2_decap_8
XFILLER_30_424 VPWR VGND sg13g2_fill_1
XFILLER_30_468 VPWR VGND sg13g2_fill_2
XFILLER_11_671 VPWR VGND sg13g2_decap_8
XFILLER_7_686 VPWR VGND sg13g2_fill_1
X_3370_ net746 _1047_ _0362_ VPWR VGND sg13g2_nor2_1
XFILLER_3_892 VPWR VGND sg13g2_decap_8
X_5040_ net164 VGND VPWR _0468_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\]
+ _0125_ sg13g2_dfrbpq_1
XFILLER_22_925 VPWR VGND sg13g2_decap_8
X_4824_ net655 net707 _0254_ VPWR VGND sg13g2_nor2_1
X_4755_ net656 net708 _0185_ VPWR VGND sg13g2_nor2_1
XFILLER_21_457 VPWR VGND sg13g2_decap_8
X_3706_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\] net566 _1375_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_30_980 VPWR VGND sg13g2_decap_8
X_4686_ net676 net728 _0116_ VPWR VGND sg13g2_nor2_1
X_3637_ _1301_ _1302_ _1304_ _1305_ _1306_ VPWR VGND sg13g2_nor4_1
X_3568_ _1222_ _1226_ _1237_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_328 VPWR VGND sg13g2_fill_2
XFILLER_0_317 VPWR VGND sg13g2_fill_1
X_3499_ _1156_ _1157_ _1164_ _1165_ _1168_ VPWR VGND sg13g2_nor4_1
X_5238_ net801 VGND VPWR net416 _0004_ clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
X_5169_ net175 VGND VPWR _0593_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\]
+ _0241_ sg13g2_dfrbpq_1
XFILLER_17_11 VPWR VGND sg13g2_fill_2
XFILLER_44_516 VPWR VGND sg13g2_fill_2
XFILLER_40_711 VPWR VGND sg13g2_fill_2
XFILLER_13_947 VPWR VGND sg13g2_decap_8
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_40_799 VPWR VGND sg13g2_fill_1
XFILLER_32_1024 VPWR VGND sg13g2_fill_1
XFILLER_3_100 VPWR VGND sg13g2_fill_1
XFILLER_4_645 VPWR VGND sg13g2_decap_8
XFILLER_3_166 VPWR VGND sg13g2_decap_8
XFILLER_0_873 VPWR VGND sg13g2_decap_8
Xhold6 serialize.n420\[1\] VPWR VGND net411 sg13g2_dlygate4sd3_1
XFILLER_48_844 VPWR VGND sg13g2_decap_8
XFILLER_47_398 VPWR VGND sg13g2_fill_2
XFILLER_16_785 VPWR VGND sg13g2_fill_2
XFILLER_43_582 VPWR VGND sg13g2_decap_8
X_2870_ net769 videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\] _0768_ _0451_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_722 VPWR VGND sg13g2_fill_2
XFILLER_31_755 VPWR VGND sg13g2_decap_8
XFILLER_31_788 VPWR VGND sg13g2_decap_4
XFILLER_8_940 VPWR VGND sg13g2_decap_8
XFILLER_30_276 VPWR VGND sg13g2_decap_8
X_4540_ _2167_ _2164_ _2169_ VPWR VGND sg13g2_xor2_1
X_4471_ _2093_ VPWR _2105_ VGND _2081_ _2092_ sg13g2_o21ai_1
X_3422_ videogen.fancy_shader.video_y\[8\] net609 _1091_ VPWR VGND sg13g2_and2_1
X_3353_ videogen.fancy_shader.video_y\[7\] videogen.fancy_shader.video_y\[6\] videogen.fancy_shader.video_y\[5\]
+ videogen.fancy_shader.video_y\[4\] _1035_ VPWR VGND sg13g2_nor4_1
X_3284_ _0975_ _0979_ _0336_ VPWR VGND sg13g2_nor2_1
X_5023_ net198 VGND VPWR _0451_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[2\]
+ _0108_ sg13g2_dfrbpq_1
XFILLER_39_855 VPWR VGND sg13g2_fill_2
XFILLER_38_343 VPWR VGND sg13g2_fill_1
X_5203__373 VPWR VGND net373 sg13g2_tiehi
XFILLER_26_549 VPWR VGND sg13g2_fill_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
X_4807_ net660 net712 _0237_ VPWR VGND sg13g2_nor2_1
X_5017__210 VPWR VGND net210 sg13g2_tiehi
X_2999_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[2\] _0802_ _0281_
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_276 VPWR VGND sg13g2_decap_4
X_4738_ net674 net726 _0168_ VPWR VGND sg13g2_nor2_1
X_4669_ net653 net705 _0099_ VPWR VGND sg13g2_nor2_1
XFILLER_1_604 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_114 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
X_4928__366 VPWR VGND net366 sg13g2_tiehi
XFILLER_29_332 VPWR VGND sg13g2_decap_4
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_17_549 VPWR VGND sg13g2_fill_2
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_9_715 VPWR VGND sg13g2_decap_4
XFILLER_13_755 VPWR VGND sg13g2_fill_2
XFILLER_13_766 VPWR VGND sg13g2_decap_8
XFILLER_8_225 VPWR VGND sg13g2_fill_1
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_0_670 VPWR VGND sg13g2_decap_8
X_4864__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_35_313 VPWR VGND sg13g2_fill_2
XFILLER_36_858 VPWR VGND sg13g2_decap_8
XFILLER_35_324 VPWR VGND sg13g2_fill_1
X_3971_ _1638_ VPWR _1639_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[0\]
+ net553 sg13g2_o21ai_1
X_2922_ _0783_ _0722_ _0781_ VPWR VGND sg13g2_nand2_2
XFILLER_16_593 VPWR VGND sg13g2_fill_2
XFILLER_31_530 VPWR VGND sg13g2_fill_2
X_2853_ _0765_ VPWR _0464_ VGND _0632_ _0764_ sg13g2_o21ai_1
X_2784_ _0737_ _0745_ _0749_ VPWR VGND sg13g2_nor2_2
X_4523_ _2153_ _2152_ _2134_ VPWR VGND sg13g2_nand2b_1
X_4454_ tmds_green.dc_balancing_reg\[2\] _2088_ _2089_ VPWR VGND sg13g2_nor2b_1
X_4898__54 VPWR VGND net54 sg13g2_tiehi
Xfanout705 net706 net705 VPWR VGND sg13g2_buf_8
X_3405_ VGND VPWR _1074_ _1073_ _1009_ sg13g2_or2_1
X_4385_ _2006_ _2027_ _2030_ VPWR VGND sg13g2_and2_1
Xfanout716 net718 net716 VPWR VGND sg13g2_buf_1
Xfanout738 net744 net738 VPWR VGND sg13g2_buf_8
X_3336_ _1024_ net795 _1023_ VPWR VGND sg13g2_nand2_1
Xfanout727 net733 net727 VPWR VGND sg13g2_buf_8
Xfanout749 net750 net749 VPWR VGND sg13g2_buf_2
X_5006_ net232 VGND VPWR _0434_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[1\]
+ _0091_ sg13g2_dfrbpq_1
XFILLER_39_652 VPWR VGND sg13g2_decap_8
X_3267_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0939_ _0969_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_22_1023 VPWR VGND sg13g2_decap_4
X_3198_ _0923_ net797 VPWR VGND _0922_ sg13g2_nand2b_2
XFILLER_35_880 VPWR VGND sg13g2_fill_1
X_4958__326 VPWR VGND net326 sg13g2_tiehi
XFILLER_14_56 VPWR VGND sg13g2_fill_2
XFILLER_10_769 VPWR VGND sg13g2_fill_1
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_39_20 VPWR VGND sg13g2_decap_8
XFILLER_18_803 VPWR VGND sg13g2_fill_2
XFILLER_29_162 VPWR VGND sg13g2_fill_2
XFILLER_44_110 VPWR VGND sg13g2_fill_2
XFILLER_32_305 VPWR VGND sg13g2_fill_2
XFILLER_44_198 VPWR VGND sg13g2_fill_1
XFILLER_13_530 VPWR VGND sg13g2_fill_2
XFILLER_40_382 VPWR VGND sg13g2_fill_1
XFILLER_45_1023 VPWR VGND sg13g2_fill_2
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_4170_ _1832_ _1816_ _1818_ VPWR VGND sg13g2_xnor2_1
X_3121_ net796 VPWR _0854_ VGND net739 net432 sg13g2_o21ai_1
XFILLER_49_994 VPWR VGND sg13g2_decap_8
X_3052_ _0839_ _0837_ _0838_ VPWR VGND sg13g2_nand2_1
XFILLER_36_644 VPWR VGND sg13g2_decap_8
XFILLER_24_817 VPWR VGND sg13g2_decap_8
X_5072__35 VPWR VGND net35 sg13g2_tiehi
X_3954_ _1622_ net593 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_32_850 VPWR VGND sg13g2_decap_8
X_2905_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[0\] net788 _0778_ _0425_
+ VPWR VGND sg13g2_mux2_1
X_3885_ net618 VPWR _1554_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[3\]
+ net561 sg13g2_o21ai_1
XFILLER_32_883 VPWR VGND sg13g2_fill_1
X_2836_ _0761_ _0722_ _0757_ VPWR VGND sg13g2_nand2_2
X_2767_ net545 _0695_ _0697_ _0744_ VPWR VGND sg13g2_nor3_2
XFILLER_2_209 VPWR VGND sg13g2_decap_8
X_2698_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\] net762 _0725_ _0588_
+ VPWR VGND sg13g2_mux2_1
X_4506_ tmds_blue.n126 tmds_blue.n132 _2136_ VPWR VGND sg13g2_and2_1
X_4437_ VGND VPWR net604 net605 _0617_ _2069_ sg13g2_a21oi_1
XFILLER_6_90 VPWR VGND sg13g2_fill_1
Xfanout546 _0691_ net546 VPWR VGND sg13g2_buf_2
Xfanout557 net560 net557 VPWR VGND sg13g2_buf_8
X_4368_ _2012_ _1996_ _2014_ VPWR VGND sg13g2_xor2_1
X_3319_ _1009_ _0999_ _1008_ VPWR VGND sg13g2_xnor2_1
X_4299_ VPWR _1961_ _1960_ VGND sg13g2_inv_1
Xfanout579 net582 net579 VPWR VGND sg13g2_buf_8
Xfanout568 net570 net568 VPWR VGND sg13g2_buf_8
XFILLER_15_828 VPWR VGND sg13g2_decap_8
XFILLER_26_154 VPWR VGND sg13g2_fill_1
XFILLER_27_666 VPWR VGND sg13g2_decap_8
XFILLER_27_677 VPWR VGND sg13g2_fill_1
XFILLER_41_135 VPWR VGND sg13g2_decap_8
XFILLER_22_382 VPWR VGND sg13g2_fill_2
XFILLER_22_393 VPWR VGND sg13g2_decap_4
XFILLER_41_98 VPWR VGND sg13g2_fill_1
XFILLER_41_87 VPWR VGND sg13g2_decap_8
XFILLER_2_710 VPWR VGND sg13g2_fill_2
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_213 VPWR VGND sg13g2_fill_2
XFILLER_46_986 VPWR VGND sg13g2_decap_8
XFILLER_18_688 VPWR VGND sg13g2_fill_1
XFILLER_40_190 VPWR VGND sg13g2_fill_2
X_3670_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\] net574 _1339_ VPWR
+ VGND sg13g2_nor2_1
X_2621_ videogen.fancy_shader.video_y\[9\] _0638_ _0673_ _0674_ VPWR VGND sg13g2_nor3_1
X_4222_ _1884_ _1139_ _1883_ VPWR VGND sg13g2_xnor2_1
X_4153_ _1812_ _1813_ _1815_ VPWR VGND sg13g2_nor2b_1
X_4948__336 VPWR VGND net336 sg13g2_tiehi
X_3104_ net422 red_tmds_par\[2\] net696 serialize.n427\[2\] VPWR VGND sg13g2_mux2_1
X_4084_ _1739_ _1742_ _1707_ _1749_ VPWR VGND sg13g2_nand3_1
X_3035_ VGND VPWR net595 net8 net549 net628 sg13g2_a21oi_2
XFILLER_37_986 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_decap_8
XFILLER_36_452 VPWR VGND sg13g2_fill_2
X_4986_ net274 VGND VPWR _0414_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\]
+ _0071_ sg13g2_dfrbpq_1
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_24_658 VPWR VGND sg13g2_decap_8
X_3937_ _1604_ VPWR _1605_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\]
+ net559 sg13g2_o21ai_1
X_3868_ net596 VPWR _1537_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\]
+ net556 sg13g2_o21ai_1
X_4955__329 VPWR VGND net329 sg13g2_tiehi
X_2819_ _0707_ _0745_ _0756_ VPWR VGND sg13g2_nor2_2
X_3799_ net612 VPWR _1468_ VGND _1463_ _1467_ sg13g2_o21ai_1
XFILLER_11_79 VPWR VGND sg13g2_decap_4
XFILLER_4_1009 VPWR VGND sg13g2_decap_8
XFILLER_19_408 VPWR VGND sg13g2_fill_2
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_43_901 VPWR VGND sg13g2_decap_4
XFILLER_28_964 VPWR VGND sg13g2_decap_8
XFILLER_43_934 VPWR VGND sg13g2_decap_8
XFILLER_42_400 VPWR VGND sg13g2_decap_8
X_4999__245 VPWR VGND net245 sg13g2_tiehi
X_5025__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_27_474 VPWR VGND sg13g2_fill_2
X_5099__295 VPWR VGND net295 sg13g2_tiehi
XFILLER_15_669 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_11_864 VPWR VGND sg13g2_fill_1
XFILLER_7_846 VPWR VGND sg13g2_fill_1
XFILLER_10_385 VPWR VGND sg13g2_fill_2
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_7 VPWR VGND sg13g2_fill_1
XFILLER_46_750 VPWR VGND sg13g2_decap_4
X_4982__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_19_986 VPWR VGND sg13g2_decap_8
X_4840_ net151 VGND VPWR _0268_ videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[1\]
+ _0007_ sg13g2_dfrbpq_1
XFILLER_34_978 VPWR VGND sg13g2_decap_8
X_4771_ net683 net734 _0201_ VPWR VGND sg13g2_nor2_1
X_3722_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[2\] net588 _1391_ VPWR
+ VGND sg13g2_nor2_1
X_3653_ _1321_ VPWR _1322_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\]
+ net580 sg13g2_o21ai_1
X_5115__229 VPWR VGND net229 sg13g2_tiehi
X_2604_ VPWR _0660_ videogen.test_lut_thingy.gol_counter_reg\[1\] VGND sg13g2_inv_1
X_3584_ _1248_ _1249_ _1252_ _1253_ VPWR VGND sg13g2_nor3_1
X_5185_ net242 VGND VPWR _0609_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[3\]
+ _0257_ sg13g2_dfrbpq_1
X_4205_ _1855_ _1853_ _1867_ VPWR VGND sg13g2_xor2_1
X_5161__238 VPWR VGND net238 sg13g2_tiehi
XFILLER_3_91 VPWR VGND sg13g2_decap_8
X_4136_ _1798_ _1697_ _1594_ VPWR VGND sg13g2_nand2b_1
XFILLER_29_706 VPWR VGND sg13g2_fill_1
XFILLER_28_227 VPWR VGND sg13g2_decap_8
X_4067_ _1731_ VPWR _1732_ VGND _1726_ _1730_ sg13g2_o21ai_1
X_3018_ videogen.fancy_shader.video_x\[4\] _0812_ _0814_ VPWR VGND sg13g2_and2_1
XFILLER_25_956 VPWR VGND sg13g2_decap_8
X_4969_ net307 VGND VPWR _0397_ videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[0\]
+ _0054_ sg13g2_dfrbpq_1
XFILLER_22_12 VPWR VGND sg13g2_fill_1
XFILLER_4_805 VPWR VGND sg13g2_fill_1
XFILLER_4_827 VPWR VGND sg13g2_decap_8
XFILLER_3_337 VPWR VGND sg13g2_decap_8
XFILLER_47_536 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_fill_2
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_43_775 VPWR VGND sg13g2_fill_1
XFILLER_42_241 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
XFILLER_15_499 VPWR VGND sg13g2_decap_8
XFILLER_11_694 VPWR VGND sg13g2_fill_1
X_4938__346 VPWR VGND net346 sg13g2_tiehi
XFILLER_3_871 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_4945__339 VPWR VGND net339 sg13g2_tiehi
XFILLER_19_761 VPWR VGND sg13g2_fill_1
XFILLER_19_772 VPWR VGND sg13g2_decap_4
XFILLER_34_720 VPWR VGND sg13g2_fill_2
XFILLER_22_904 VPWR VGND sg13g2_decap_8
X_4823_ net652 net704 _0253_ VPWR VGND sg13g2_nor2_1
X_4754_ net673 net708 _0184_ VPWR VGND sg13g2_nor2_1
X_3705_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\] net588 _1374_ VPWR
+ VGND sg13g2_nor2_1
X_4685_ net679 net731 _0115_ VPWR VGND sg13g2_nor2_1
X_3636_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\] net573 _1305_ VPWR
+ VGND sg13g2_nor2_1
X_3567_ _1233_ _1234_ _1236_ VPWR VGND sg13g2_and2_1
X_5237_ net801 VGND VPWR serialize.n433\[1\] serialize.bit_cnt\[1\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3498_ _1164_ _1165_ _1167_ VPWR VGND sg13g2_nor2_1
XFILLER_29_514 VPWR VGND sg13g2_fill_1
X_5168_ net183 VGND VPWR _0592_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\]
+ _0240_ sg13g2_dfrbpq_1
X_5099_ net295 VGND VPWR _0523_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[1\]
+ _0171_ sg13g2_dfrbpq_1
X_4119_ _1778_ _1780_ _1236_ _1784_ VPWR VGND _1781_ sg13g2_nand4_1
XFILLER_25_753 VPWR VGND sg13g2_fill_1
XFILLER_40_701 VPWR VGND sg13g2_fill_1
XFILLER_13_926 VPWR VGND sg13g2_decap_8
XFILLER_12_436 VPWR VGND sg13g2_fill_2
XFILLER_8_418 VPWR VGND sg13g2_decap_4
XFILLER_21_992 VPWR VGND sg13g2_decap_8
XFILLER_4_635 VPWR VGND sg13g2_fill_1
XFILLER_0_852 VPWR VGND sg13g2_decap_8
XFILLER_48_823 VPWR VGND sg13g2_decap_8
Xhold7 serialize.bit_cnt\[0\] VPWR VGND net412 sg13g2_dlygate4sd3_1
XFILLER_35_506 VPWR VGND sg13g2_fill_1
XFILLER_28_580 VPWR VGND sg13g2_decap_8
XFILLER_28_591 VPWR VGND sg13g2_fill_2
XFILLER_43_594 VPWR VGND sg13g2_decap_4
XFILLER_15_274 VPWR VGND sg13g2_fill_2
X_4470_ _2104_ _2102_ _2103_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_996 VPWR VGND sg13g2_decap_8
XFILLER_7_484 VPWR VGND sg13g2_fill_2
X_3421_ VPWR _1090_ net544 VGND sg13g2_inv_1
X_3352_ _1032_ _1034_ _0357_ VPWR VGND sg13g2_nor2_1
X_3283_ _0979_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] _0977_ VPWR
+ VGND sg13g2_xnor2_1
XFILLER_39_845 VPWR VGND sg13g2_decap_4
X_5022_ net200 VGND VPWR _0450_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[1\]
+ _0107_ sg13g2_dfrbpq_1
XFILLER_19_580 VPWR VGND sg13g2_decap_8
X_4806_ net653 net705 _0236_ VPWR VGND sg13g2_nor2_1
X_2998_ net754 videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[3\] _0802_ _0282_
+ VPWR VGND sg13g2_mux2_1
X_4737_ net677 net729 _0167_ VPWR VGND sg13g2_nor2_1
X_4668_ net653 net705 _0098_ VPWR VGND sg13g2_nor2_1
X_3619_ _1235_ _1275_ _1288_ VPWR VGND sg13g2_nor2_1
X_4599_ net661 net713 _0029_ VPWR VGND sg13g2_nor2_1
XFILLER_0_126 VPWR VGND sg13g2_decap_4
XFILLER_29_311 VPWR VGND sg13g2_fill_1
XFILLER_44_347 VPWR VGND sg13g2_fill_1
XFILLER_12_222 VPWR VGND sg13g2_decap_8
XFILLER_40_575 VPWR VGND sg13g2_fill_2
XFILLER_8_237 VPWR VGND sg13g2_decap_4
XFILLER_12_255 VPWR VGND sg13g2_decap_8
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_5_37 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_4
XFILLER_47_141 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
X_3970_ _1638_ net594 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_43_380 VPWR VGND sg13g2_decap_4
X_2921_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\] _0782_ _0413_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_542 VPWR VGND sg13g2_fill_2
XFILLER_31_553 VPWR VGND sg13g2_decap_8
X_2852_ _0765_ net757 _0764_ VPWR VGND sg13g2_nand2_1
X_2783_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[0\] net790 _0748_ _0526_
+ VPWR VGND sg13g2_mux2_1
X_4522_ _2152_ _2142_ _2150_ VPWR VGND sg13g2_xnor2_1
X_4453_ _2088_ _2086_ VPWR VGND _2084_ sg13g2_nand2b_2
X_3404_ _1073_ _1071_ _1072_ VPWR VGND sg13g2_nand2_2
X_4901__48 VPWR VGND net48 sg13g2_tiehi
Xfanout706 net724 net706 VPWR VGND sg13g2_buf_2
X_4384_ _2029_ _2007_ _2028_ VPWR VGND sg13g2_nand2_1
Xfanout717 net718 net717 VPWR VGND sg13g2_buf_8
X_3335_ videogen.fancy_shader.n646\[5\] _1019_ videogen.fancy_shader.n646\[6\] _1023_
+ VPWR VGND sg13g2_nand3_1
Xfanout728 net733 net728 VPWR VGND sg13g2_buf_1
Xfanout739 net740 net739 VPWR VGND sg13g2_buf_8
X_3266_ _0939_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0968_ VPWR
+ VGND sg13g2_nor2b_1
X_5005_ net234 VGND VPWR _0433_ videogen.test_lut_thingy.pixel_feeder_inst.row\[51\]\[0\]
+ _0090_ sg13g2_dfrbpq_1
XFILLER_22_1002 VPWR VGND sg13g2_decap_8
XFILLER_38_152 VPWR VGND sg13g2_fill_1
XFILLER_38_141 VPWR VGND sg13g2_decap_8
X_3197_ _0922_ _0806_ _0814_ _0921_ VPWR VGND sg13g2_and3_2
XFILLER_14_35 VPWR VGND sg13g2_decap_8
XFILLER_34_380 VPWR VGND sg13g2_fill_1
XFILLER_10_704 VPWR VGND sg13g2_fill_1
XFILLER_14_79 VPWR VGND sg13g2_decap_8
X_5145__37 VPWR VGND net37 sg13g2_tiehi
XFILLER_2_936 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_39_76 VPWR VGND sg13g2_fill_1
XFILLER_17_303 VPWR VGND sg13g2_decap_8
XFILLER_45_645 VPWR VGND sg13g2_decap_4
XFILLER_18_837 VPWR VGND sg13g2_fill_2
XFILLER_44_144 VPWR VGND sg13g2_decap_4
XFILLER_17_369 VPWR VGND sg13g2_decap_8
XFILLER_26_881 VPWR VGND sg13g2_decap_8
XFILLER_41_862 VPWR VGND sg13g2_fill_2
XFILLER_13_542 VPWR VGND sg13g2_fill_2
XFILLER_9_513 VPWR VGND sg13g2_fill_1
XFILLER_13_586 VPWR VGND sg13g2_decap_4
XFILLER_9_546 VPWR VGND sg13g2_fill_1
X_5035__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_5_785 VPWR VGND sg13g2_fill_2
X_3120_ tmds_blue.dc_balancing_reg\[0\] _0852_ _0264_ VPWR VGND sg13g2_and2_1
XFILLER_1_991 VPWR VGND sg13g2_decap_8
XFILLER_49_973 VPWR VGND sg13g2_decap_8
X_3051_ _0694_ net549 videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0838_
+ VPWR VGND sg13g2_a21o_1
X_3953_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\] net550 _1621_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_16_380 VPWR VGND sg13g2_decap_8
X_2904_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[1\] net777 _0778_ _0426_
+ VPWR VGND sg13g2_mux2_1
X_3884_ net614 _1547_ _1552_ _1553_ VPWR VGND sg13g2_nor3_1
X_2835_ net784 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[0\] _0760_ _0477_
+ VPWR VGND sg13g2_mux2_1
X_2766_ _0695_ _0697_ _0743_ VPWR VGND sg13g2_nor2_2
X_2697_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\] net754 _0725_ _0589_
+ VPWR VGND sg13g2_mux2_1
X_4505_ net572 _2135_ _0624_ VPWR VGND sg13g2_nor2_1
X_4436_ VGND VPWR net605 _2074_ _0616_ _2064_ sg13g2_a21oi_1
X_4367_ _1996_ _2012_ _2013_ VPWR VGND sg13g2_nor2_1
X_3318_ VGND VPWR _1008_ _1007_ _1000_ sg13g2_or2_1
Xfanout547 _0881_ net547 VPWR VGND sg13g2_buf_8
X_4298_ _1942_ _1943_ _1955_ _1959_ _1960_ VPWR VGND sg13g2_and4_1
Xfanout558 net560 net558 VPWR VGND sg13g2_buf_8
Xfanout569 net570 net569 VPWR VGND sg13g2_buf_8
X_3249_ VPWR _0957_ _0956_ VGND sg13g2_inv_1
XFILLER_26_111 VPWR VGND sg13g2_fill_2
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_15_818 VPWR VGND sg13g2_fill_2
XFILLER_41_103 VPWR VGND sg13g2_decap_4
XFILLER_26_188 VPWR VGND sg13g2_decap_8
XFILLER_42_648 VPWR VGND sg13g2_decap_8
XFILLER_41_125 VPWR VGND sg13g2_decap_4
XFILLER_22_361 VPWR VGND sg13g2_fill_1
XFILLER_10_512 VPWR VGND sg13g2_fill_1
XFILLER_23_895 VPWR VGND sg13g2_decap_8
XFILLER_41_66 VPWR VGND sg13g2_decap_4
XFILLER_41_55 VPWR VGND sg13g2_decap_8
XFILLER_10_567 VPWR VGND sg13g2_decap_8
XFILLER_9_2 VPWR VGND sg13g2_fill_1
XFILLER_49_269 VPWR VGND sg13g2_fill_2
XFILLER_46_965 VPWR VGND sg13g2_decap_8
XFILLER_17_144 VPWR VGND sg13g2_decap_4
XFILLER_17_155 VPWR VGND sg13g2_fill_1
XFILLER_45_486 VPWR VGND sg13g2_fill_2
XFILLER_14_862 VPWR VGND sg13g2_fill_2
XFILLER_13_372 VPWR VGND sg13g2_decap_8
XFILLER_9_376 VPWR VGND sg13g2_decap_8
X_2620_ videogen.fancy_shader.video_y\[6\] videogen.fancy_shader.video_y\[5\] videogen.fancy_shader.video_y\[7\]
+ _0673_ VPWR VGND sg13g2_nand3_1
XFILLER_5_571 VPWR VGND sg13g2_decap_8
X_4221_ _1883_ _1809_ _1882_ VPWR VGND sg13g2_xnor2_1
X_4152_ _1810_ _1813_ _1808_ _1814_ VPWR VGND sg13g2_nand3_1
X_3103_ net441 red_tmds_par\[1\] net699 serialize.n427\[1\] VPWR VGND sg13g2_mux2_1
X_4083_ _1736_ _1728_ _1748_ VPWR VGND sg13g2_xor2_1
X_3034_ serialize.bit_cnt\[1\] net412 net415 serialize.n410 VPWR VGND sg13g2_nor3_1
XFILLER_24_626 VPWR VGND sg13g2_decap_8
XFILLER_36_475 VPWR VGND sg13g2_decap_4
X_4985_ net276 VGND VPWR _0413_ videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[0\]
+ _0070_ sg13g2_dfrbpq_1
XFILLER_23_169 VPWR VGND sg13g2_decap_8
X_3936_ _1604_ net594 videogen.test_lut_thingy.pixel_feeder_inst.row\[16\]\[0\] VPWR
+ VGND sg13g2_nand2b_1
X_3867_ videogen.test_lut_thingy.pixel_feeder_inst.row\[32\]\[3\] net585 _1536_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_31_180 VPWR VGND sg13g2_decap_4
X_2818_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[0\] net786 _0755_ _0489_
+ VPWR VGND sg13g2_mux2_1
X_3798_ net615 VPWR _1467_ VGND _1464_ _1466_ sg13g2_o21ai_1
XFILLER_3_508 VPWR VGND sg13g2_decap_8
X_2749_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\] net781 _0739_ _0551_
+ VPWR VGND sg13g2_mux2_1
X_4419_ _2062_ net602 _2060_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_943 VPWR VGND sg13g2_decap_8
XFILLER_15_615 VPWR VGND sg13g2_fill_2
XFILLER_36_88 VPWR VGND sg13g2_fill_1
XFILLER_36_99 VPWR VGND sg13g2_decap_8
XFILLER_14_158 VPWR VGND sg13g2_fill_1
XFILLER_23_692 VPWR VGND sg13g2_fill_1
XFILLER_6_335 VPWR VGND sg13g2_fill_2
XFILLER_2_574 VPWR VGND sg13g2_decap_4
XFILLER_18_420 VPWR VGND sg13g2_fill_1
XFILLER_19_965 VPWR VGND sg13g2_decap_8
X_5004__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_34_957 VPWR VGND sg13g2_decap_8
XFILLER_20_117 VPWR VGND sg13g2_fill_1
X_4770_ net683 net734 _0200_ VPWR VGND sg13g2_nor2_1
X_3721_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[2\] net573 _1390_ VPWR
+ VGND sg13g2_nor2_1
X_3652_ _1319_ _1320_ _1321_ VPWR VGND sg13g2_nor2_1
X_4954__330 VPWR VGND net330 sg13g2_tiehi
X_2603_ _0659_ videogen.test_lut_thingy.pixel_feeder_inst.state\[2\] VPWR VGND sg13g2_inv_2
X_3583_ _1252_ net544 _1251_ VPWR VGND sg13g2_nand2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5184_ net258 VGND VPWR _0608_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[2\]
+ _0256_ sg13g2_dfrbpq_1
X_4204_ VGND VPWR _1853_ _1864_ _1866_ _1861_ sg13g2_a21oi_1
X_4135_ _0378_ _1790_ _1797_ VPWR VGND sg13g2_nand2_2
X_4961__323 VPWR VGND net323 sg13g2_tiehi
X_4066_ _1731_ _1719_ _1723_ VPWR VGND sg13g2_nand2_1
X_3017_ _0813_ videogen.fancy_shader.video_x\[3\] _0811_ VPWR VGND sg13g2_nand2_1
XFILLER_25_935 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_40_905 VPWR VGND sg13g2_fill_2
XFILLER_24_489 VPWR VGND sg13g2_decap_4
X_4968_ net309 VGND VPWR _0396_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\]
+ _0053_ sg13g2_dfrbpq_1
X_4899_ net52 VGND VPWR _0327_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[3\]
+ net630 sg13g2_dfrbpq_2
X_3919_ _0644_ _1576_ _1587_ _1588_ VPWR VGND sg13g2_nor3_1
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_32 VPWR VGND sg13g2_fill_1
XFILLER_28_740 VPWR VGND sg13g2_fill_1
XFILLER_16_924 VPWR VGND sg13g2_decap_8
XFILLER_28_762 VPWR VGND sg13g2_fill_2
XFILLER_28_773 VPWR VGND sg13g2_decap_4
XFILLER_43_732 VPWR VGND sg13g2_fill_1
XFILLER_15_478 VPWR VGND sg13g2_decap_4
XFILLER_24_990 VPWR VGND sg13g2_decap_8
XFILLER_30_415 VPWR VGND sg13g2_decap_8
XFILLER_31_949 VPWR VGND sg13g2_decap_8
XFILLER_7_633 VPWR VGND sg13g2_fill_2
XFILLER_10_150 VPWR VGND sg13g2_fill_1
XFILLER_10_172 VPWR VGND sg13g2_fill_1
XFILLER_6_176 VPWR VGND sg13g2_decap_4
XFILLER_6_198 VPWR VGND sg13g2_decap_4
XFILLER_3_850 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_fill_1
XFILLER_46_570 VPWR VGND sg13g2_decap_8
X_4822_ net654 net706 _0252_ VPWR VGND sg13g2_nor2_1
XFILLER_21_426 VPWR VGND sg13g2_decap_4
X_4753_ net673 net725 _0183_ VPWR VGND sg13g2_nor2_1
X_3704_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\] net556 _1373_ VPWR
+ VGND sg13g2_nor2_1
X_4684_ net681 net728 _0114_ VPWR VGND sg13g2_nor2_1
X_3635_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[2\] net567 _1304_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_1_809 VPWR VGND sg13g2_decap_8
X_3566_ _1235_ _1233_ _1234_ VPWR VGND sg13g2_nand2_2
X_3497_ VGND VPWR _1166_ _1165_ _1164_ sg13g2_or2_1
X_5236_ net801 VGND VPWR serialize.n433\[0\] serialize.bit_cnt\[0\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_2
X_5167_ net191 VGND VPWR _0591_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\]
+ _0239_ sg13g2_dfrbpq_1
X_5098_ net299 VGND VPWR _0522_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[0\]
+ _0170_ sg13g2_dfrbpq_1
X_4118_ _1778_ _1782_ _1783_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_518 VPWR VGND sg13g2_fill_1
X_4049_ _1145_ _1709_ _1714_ VPWR VGND sg13g2_and2_1
XFILLER_17_79 VPWR VGND sg13g2_decap_8
XFILLER_13_905 VPWR VGND sg13g2_decap_8
XFILLER_40_713 VPWR VGND sg13g2_fill_1
X_5172__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_24_297 VPWR VGND sg13g2_decap_4
XFILLER_21_971 VPWR VGND sg13g2_decap_8
XFILLER_4_614 VPWR VGND sg13g2_decap_8
XFILLER_0_831 VPWR VGND sg13g2_decap_8
Xhold8 serialize.n420\[4\] VPWR VGND net413 sg13g2_dlygate4sd3_1
XFILLER_48_879 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_fill_2
X_4944__340 VPWR VGND net340 sg13g2_tiehi
XFILLER_35_529 VPWR VGND sg13g2_decap_4
XFILLER_43_562 VPWR VGND sg13g2_decap_8
XFILLER_16_787 VPWR VGND sg13g2_fill_1
XFILLER_31_746 VPWR VGND sg13g2_fill_2
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_8_975 VPWR VGND sg13g2_decap_8
XFILLER_7_496 VPWR VGND sg13g2_decap_8
X_3420_ _1088_ _1082_ _1089_ VPWR VGND sg13g2_xor2_1
X_4951__333 VPWR VGND net333 sg13g2_tiehi
X_3351_ net798 VPWR _1034_ VGND videogen.fancy_shader.video_y\[1\] _1030_ sg13g2_o21ai_1
XFILLER_3_691 VPWR VGND sg13g2_decap_8
X_3282_ _0975_ _0977_ _0978_ _0335_ VPWR VGND sg13g2_nor3_1
X_5021_ net202 VGND VPWR _0449_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\]
+ _0106_ sg13g2_dfrbpq_1
XFILLER_39_857 VPWR VGND sg13g2_fill_1
XFILLER_0_60 VPWR VGND sg13g2_decap_8
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_decap_4
X_4805_ net660 net712 _0235_ VPWR VGND sg13g2_nor2_1
X_2997_ _0802_ _0781_ VPWR VGND _0737_ sg13g2_nand2b_2
X_4736_ net678 net732 _0166_ VPWR VGND sg13g2_nor2_1
X_4667_ net685 net737 _0097_ VPWR VGND sg13g2_nor2_1
X_3618_ _1284_ _1285_ _1286_ _1287_ VPWR VGND sg13g2_nor3_1
X_4598_ net662 net714 _0028_ VPWR VGND sg13g2_nor2_1
XFILLER_0_105 VPWR VGND sg13g2_fill_1
X_3549_ VGND VPWR _1211_ _1215_ _1218_ _1217_ sg13g2_a21oi_1
X_5219_ net803 VGND VPWR serialize.n431\[1\] serialize.n461 clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_34 VPWR VGND sg13g2_decap_8
XFILLER_45_816 VPWR VGND sg13g2_decap_4
XFILLER_38_890 VPWR VGND sg13g2_fill_1
XFILLER_12_201 VPWR VGND sg13g2_decap_8
XFILLER_40_532 VPWR VGND sg13g2_decap_8
XFILLER_8_205 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_12_289 VPWR VGND sg13g2_decap_4
XFILLER_5_923 VPWR VGND sg13g2_decap_8
X_5111__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_10_8 VPWR VGND sg13g2_decap_8
XFILLER_36_805 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_fill_1
X_2920_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\] _0782_ _0414_
+ VPWR VGND sg13g2_mux2_1
X_4979__288 VPWR VGND net288 sg13g2_tiehi
XFILLER_31_521 VPWR VGND sg13g2_decap_4
XFILLER_31_532 VPWR VGND sg13g2_fill_1
XFILLER_15_1010 VPWR VGND sg13g2_decap_8
X_2851_ _0726_ _0758_ _0764_ VPWR VGND sg13g2_nor2_2
X_2782_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[1\] net779 _0748_ _0527_
+ VPWR VGND sg13g2_mux2_1
X_4521_ _2151_ _2150_ _2142_ VPWR VGND sg13g2_nand2b_1
X_4452_ net601 _2083_ _2087_ VPWR VGND sg13g2_nor2_1
X_3403_ _1070_ VPWR _1072_ VGND _1067_ _1068_ sg13g2_o21ai_1
X_4383_ _2027_ _2022_ _2028_ VPWR VGND sg13g2_xor2_1
X_3334_ VGND VPWR videogen.fancy_shader.n646\[5\] _1019_ _1022_ videogen.fancy_shader.n646\[6\]
+ sg13g2_a21oi_1
Xfanout707 net708 net707 VPWR VGND sg13g2_buf_8
Xfanout729 net732 net729 VPWR VGND sg13g2_buf_8
Xfanout718 net724 net718 VPWR VGND sg13g2_buf_8
X_3265_ VGND VPWR _0967_ _0943_ _0940_ sg13g2_or2_1
X_5004_ net235 VGND VPWR _0432_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[3\]
+ _0089_ sg13g2_dfrbpq_1
X_3196_ net629 videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\]
+ _0921_ VPWR VGND sg13g2_nor3_1
XFILLER_38_197 VPWR VGND sg13g2_fill_1
XFILLER_38_186 VPWR VGND sg13g2_fill_2
XFILLER_14_58 VPWR VGND sg13g2_fill_1
X_4719_ net662 net714 _0149_ VPWR VGND sg13g2_nor2_1
XFILLER_2_915 VPWR VGND sg13g2_decap_8
XFILLER_1_425 VPWR VGND sg13g2_decap_4
XFILLER_49_418 VPWR VGND sg13g2_decap_8
XFILLER_39_55 VPWR VGND sg13g2_fill_2
XFILLER_17_348 VPWR VGND sg13g2_fill_2
X_4941__343 VPWR VGND net343 sg13g2_tiehi
XFILLER_26_860 VPWR VGND sg13g2_decap_8
XFILLER_38_1021 VPWR VGND sg13g2_decap_8
XFILLER_32_307 VPWR VGND sg13g2_fill_1
XFILLER_41_841 VPWR VGND sg13g2_decap_8
XFILLER_5_764 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_4
XFILLER_1_970 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_decap_8
X_3050_ net549 _0694_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0837_
+ VPWR VGND sg13g2_nand3_1
XFILLER_36_613 VPWR VGND sg13g2_decap_8
XFILLER_17_860 VPWR VGND sg13g2_decap_8
XFILLER_17_871 VPWR VGND sg13g2_fill_1
X_3952_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[0\] net574 _1620_ VPWR
+ VGND sg13g2_nor2_1
X_2903_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[2\] net765 _0778_ _0427_
+ VPWR VGND sg13g2_mux2_1
X_3883_ net621 _1548_ _1549_ _1551_ _1552_ VPWR VGND sg13g2_nor4_1
XFILLER_32_874 VPWR VGND sg13g2_decap_8
X_5118__217 VPWR VGND net217 sg13g2_tiehi
X_5192__179 VPWR VGND net179 sg13g2_tiehi
X_2834_ net773 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[1\] _0760_ _0478_
+ VPWR VGND sg13g2_mux2_1
X_2765_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[0\] _0742_ _0538_
+ VPWR VGND sg13g2_mux2_1
X_4504_ _2134_ _2063_ _2135_ VPWR VGND sg13g2_xor2_1
X_2696_ _0714_ _0722_ _0725_ VPWR VGND sg13g2_nor2b_2
X_4435_ _2074_ _2072_ _2073_ VPWR VGND sg13g2_xnor2_1
X_4366_ _2011_ _1999_ _2012_ VPWR VGND sg13g2_xor2_1
X_3317_ VPWR VGND _1006_ _1001_ _1002_ videogen.fancy_shader.n646\[3\] _1007_ videogen.fancy_shader.video_x\[3\]
+ sg13g2_a221oi_1
X_5164__215 VPWR VGND net215 sg13g2_tiehi
Xfanout548 _0881_ net548 VPWR VGND sg13g2_buf_1
X_4297_ _1959_ _1944_ _1954_ VPWR VGND sg13g2_nand2_1
Xfanout559 net560 net559 VPWR VGND sg13g2_buf_8
XFILLER_39_462 VPWR VGND sg13g2_fill_1
X_3248_ _0807_ _0955_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[3\] _0956_
+ VPWR VGND sg13g2_nand3_1
X_4847__141 VPWR VGND net141 sg13g2_tiehi
X_3179_ _0908_ _0907_ _0902_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_35 VPWR VGND sg13g2_fill_2
X_5101__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_22_384 VPWR VGND sg13g2_fill_1
X_4971__303 VPWR VGND net303 sg13g2_tiehi
XFILLER_2_701 VPWR VGND sg13g2_decap_4
XFILLER_2_789 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_49_215 VPWR VGND sg13g2_fill_1
XFILLER_49_259 VPWR VGND sg13g2_fill_2
XFILLER_46_944 VPWR VGND sg13g2_decap_8
XFILLER_33_627 VPWR VGND sg13g2_decap_4
XFILLER_45_498 VPWR VGND sg13g2_fill_1
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_33_649 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_4
XFILLER_13_395 VPWR VGND sg13g2_decap_8
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_4220_ VGND VPWR _1161_ _1162_ _1882_ _1879_ sg13g2_a21oi_1
X_4151_ _1803_ _1717_ _1813_ VPWR VGND sg13g2_xor2_1
X_3102_ net421 red_tmds_par\[0\] net699 serialize.n427\[0\] VPWR VGND sg13g2_mux2_1
X_4876__92 VPWR VGND net92 sg13g2_tiehi
X_4082_ VGND VPWR _1747_ _1746_ _1745_ sg13g2_or2_1
XFILLER_37_922 VPWR VGND sg13g2_decap_8
X_3033_ VGND VPWR _0659_ _0827_ _0003_ net746 sg13g2_a21oi_1
XFILLER_23_104 VPWR VGND sg13g2_fill_1
XFILLER_24_605 VPWR VGND sg13g2_decap_8
X_4984_ net278 VGND VPWR _0412_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[3\]
+ _0069_ sg13g2_dfrbpq_1
X_3935_ videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\] net569 _1603_ VPWR
+ VGND sg13g2_nor2_1
X_3866_ videogen.test_lut_thingy.pixel_feeder_inst.row\[35\]\[3\] net573 _1535_ VPWR
+ VGND sg13g2_nor2_1
X_2817_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[1\] net775 _0755_ _0490_
+ VPWR VGND sg13g2_mux2_1
X_3797_ _1465_ VPWR _1466_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\]
+ net553 sg13g2_o21ai_1
X_2748_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\] net770 _0739_ _0552_
+ VPWR VGND sg13g2_mux2_1
X_4418_ _2061_ _2058_ _2059_ VPWR VGND sg13g2_nand2_2
X_2679_ _0720_ _0646_ _0704_ _0706_ VPWR VGND sg13g2_and3_2
XFILLER_28_1020 VPWR VGND sg13g2_decap_8
X_4349_ _1996_ tmds_red.n114 _1995_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_922 VPWR VGND sg13g2_decap_8
XFILLER_14_104 VPWR VGND sg13g2_decap_8
XFILLER_27_465 VPWR VGND sg13g2_decap_4
XFILLER_28_999 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_4
XFILLER_43_969 VPWR VGND sg13g2_decap_8
XFILLER_42_468 VPWR VGND sg13g2_fill_2
XFILLER_42_457 VPWR VGND sg13g2_decap_8
XFILLER_11_800 VPWR VGND sg13g2_fill_1
XFILLER_10_310 VPWR VGND sg13g2_decap_8
XFILLER_10_321 VPWR VGND sg13g2_fill_1
XFILLER_10_354 VPWR VGND sg13g2_fill_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
X_4910__404 VPWR VGND net404 sg13g2_tiehi
XFILLER_2_553 VPWR VGND sg13g2_decap_8
XFILLER_2_597 VPWR VGND sg13g2_decap_8
X_4873__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_19_944 VPWR VGND sg13g2_decap_8
XFILLER_18_465 VPWR VGND sg13g2_fill_2
XFILLER_34_936 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_fill_2
XFILLER_42_980 VPWR VGND sg13g2_decap_8
X_3720_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[2\] net567 _1389_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_13_170 VPWR VGND sg13g2_decap_8
X_3651_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[2\] net558 _1320_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_9_196 VPWR VGND sg13g2_fill_2
X_3582_ VGND VPWR _1139_ _1166_ _1251_ _1158_ sg13g2_a21oi_1
X_2602_ VPWR _0658_ net796 VGND sg13g2_inv_1
X_5183_ net277 VGND VPWR _0607_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\]
+ _0255_ sg13g2_dfrbpq_1
X_4203_ _1864_ _1862_ _1860_ _1865_ VPWR VGND sg13g2_a21o_1
X_4134_ _1795_ _1796_ _1592_ _1797_ VPWR VGND sg13g2_nand3_1
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
XFILLER_28_218 VPWR VGND sg13g2_decap_4
XFILLER_49_590 VPWR VGND sg13g2_decap_8
X_4065_ _1717_ _1725_ _1727_ _1729_ _1730_ VPWR VGND sg13g2_and4_1
X_4844__144 VPWR VGND net144 sg13g2_tiehi
X_3016_ videogen.fancy_shader.video_x\[3\] _0811_ _0812_ VPWR VGND sg13g2_and2_1
XFILLER_25_914 VPWR VGND sg13g2_decap_8
XFILLER_36_240 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_40_928 VPWR VGND sg13g2_fill_1
XFILLER_24_479 VPWR VGND sg13g2_decap_4
X_4967_ net311 VGND VPWR _0395_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[2\]
+ _0052_ sg13g2_dfrbpq_1
XFILLER_33_980 VPWR VGND sg13g2_decap_8
X_4898_ net54 VGND VPWR _0326_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[2\]
+ net630 sg13g2_dfrbpq_2
X_3918_ net597 _1581_ _1586_ _1587_ VPWR VGND sg13g2_nor3_1
X_3849_ net612 VPWR _1518_ VGND _1512_ _1517_ sg13g2_o21ai_1
XFILLER_22_47 VPWR VGND sg13g2_decap_8
XFILLER_22_58 VPWR VGND sg13g2_decap_4
X_4851__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_44 VPWR VGND sg13g2_decap_8
X_5107__260 VPWR VGND net260 sg13g2_tiehi
XFILLER_16_903 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_decap_4
XFILLER_42_210 VPWR VGND sg13g2_fill_1
XFILLER_27_273 VPWR VGND sg13g2_fill_2
XFILLER_31_928 VPWR VGND sg13g2_decap_8
XFILLER_7_601 VPWR VGND sg13g2_fill_1
XFILLER_11_663 VPWR VGND sg13g2_fill_2
XFILLER_11_685 VPWR VGND sg13g2_decap_8
XFILLER_33_210 VPWR VGND sg13g2_fill_1
XFILLER_34_733 VPWR VGND sg13g2_decap_8
X_4821_ net653 net705 _0251_ VPWR VGND sg13g2_nor2_1
XFILLER_22_939 VPWR VGND sg13g2_decap_8
X_4752_ net673 net725 _0182_ VPWR VGND sg13g2_nor2_1
X_3703_ net596 VPWR _1372_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[39\]\[2\]
+ net578 sg13g2_o21ai_1
X_4683_ net675 net727 _0113_ VPWR VGND sg13g2_nor2_1
X_3634_ _1303_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[0\] VPWR VGND videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\]
+ sg13g2_nand2b_2
XFILLER_30_994 VPWR VGND sg13g2_decap_8
X_3565_ _1234_ videogen.fancy_shader.video_y\[0\] videogen.fancy_shader.video_x\[0\]
+ VPWR VGND sg13g2_nand2_1
X_3496_ _1127_ _1159_ _1161_ _1162_ _1165_ VPWR VGND sg13g2_and4_1
X_5235_ net799 VGND VPWR serialize.n429\[9\] serialize.n417\[7\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
X_5166_ net199 VGND VPWR _0590_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\]
+ _0238_ sg13g2_dfrbpq_1
X_5097_ net302 VGND VPWR _0521_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[3\]
+ _0169_ sg13g2_dfrbpq_1
X_4117_ _1780_ _1781_ _1236_ _1782_ VPWR VGND sg13g2_nand3_1
X_4048_ _1713_ _1711_ _1712_ VPWR VGND sg13g2_nand2_1
XFILLER_17_25 VPWR VGND sg13g2_decap_8
XFILLER_25_700 VPWR VGND sg13g2_fill_2
XFILLER_17_69 VPWR VGND sg13g2_fill_1
XFILLER_25_766 VPWR VGND sg13g2_decap_8
XFILLER_25_777 VPWR VGND sg13g2_fill_1
XFILLER_12_449 VPWR VGND sg13g2_fill_2
XFILLER_21_950 VPWR VGND sg13g2_decap_8
XFILLER_4_659 VPWR VGND sg13g2_decap_4
XFILLER_3_125 VPWR VGND sg13g2_decap_8
XFILLER_0_810 VPWR VGND sg13g2_decap_8
Xhold9 serialize.n414\[1\] VPWR VGND net414 sg13g2_dlygate4sd3_1
XFILLER_0_887 VPWR VGND sg13g2_decap_8
XFILLER_48_858 VPWR VGND sg13g2_decap_8
XFILLER_47_335 VPWR VGND sg13g2_fill_1
XFILLER_16_711 VPWR VGND sg13g2_decap_8
XFILLER_16_733 VPWR VGND sg13g2_fill_2
XFILLER_43_541 VPWR VGND sg13g2_decap_8
XFILLER_15_276 VPWR VGND sg13g2_fill_1
XFILLER_31_769 VPWR VGND sg13g2_fill_2
XFILLER_11_460 VPWR VGND sg13g2_decap_8
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_30_257 VPWR VGND sg13g2_decap_4
XFILLER_8_954 VPWR VGND sg13g2_decap_8
XFILLER_11_471 VPWR VGND sg13g2_fill_1
XFILLER_7_464 VPWR VGND sg13g2_decap_8
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
X_3350_ _1033_ _0922_ _0831_ VPWR VGND sg13g2_nand2b_1
X_5020_ net204 VGND VPWR _0448_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[3\]
+ _0105_ sg13g2_dfrbpq_1
X_3281_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\] _0818_ _0978_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_38_335 VPWR VGND sg13g2_fill_1
XFILLER_46_390 VPWR VGND sg13g2_decap_4
XFILLER_0_94 VPWR VGND sg13g2_decap_8
XFILLER_10_909 VPWR VGND sg13g2_decap_8
XFILLER_22_747 VPWR VGND sg13g2_decap_4
X_4804_ net660 net712 _0234_ VPWR VGND sg13g2_nor2_1
XFILLER_34_596 VPWR VGND sg13g2_fill_2
X_4735_ net677 net729 _0165_ VPWR VGND sg13g2_nor2_1
X_2996_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[0\] net785 _0801_ _0283_
+ VPWR VGND sg13g2_mux2_1
X_4666_ net685 net736 _0096_ VPWR VGND sg13g2_nor2_1
X_5132__161 VPWR VGND net161 sg13g2_tiehi
X_3617_ _1286_ _1236_ _1282_ VPWR VGND sg13g2_nand2_1
X_4597_ net661 net713 _0027_ VPWR VGND sg13g2_nor2_1
X_3548_ _1216_ VPWR _1217_ VGND _1198_ _1205_ sg13g2_o21ai_1
XFILLER_1_629 VPWR VGND sg13g2_fill_1
X_3479_ VGND VPWR _1147_ _1148_ _1137_ _1135_ sg13g2_a21oi_2
XFILLER_0_139 VPWR VGND sg13g2_fill_2
X_5218_ net803 VGND VPWR serialize.n431\[0\] serialize.n459 clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5149_ net377 VGND VPWR _0573_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[3\]
+ _0221_ sg13g2_dfrbpq_1
XFILLER_28_57 VPWR VGND sg13g2_fill_2
XFILLER_28_68 VPWR VGND sg13g2_decap_8
XFILLER_28_79 VPWR VGND sg13g2_fill_1
XFILLER_25_552 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_decap_8
XFILLER_13_714 VPWR VGND sg13g2_decap_8
X_5178__397 VPWR VGND net397 sg13g2_tiehi
XFILLER_40_588 VPWR VGND sg13g2_decap_8
XFILLER_12_268 VPWR VGND sg13g2_decap_8
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_4_489 VPWR VGND sg13g2_decap_8
XFILLER_47_121 VPWR VGND sg13g2_decap_4
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_48_666 VPWR VGND sg13g2_decap_8
X_2850_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[0\] net789 _0763_ _0465_
+ VPWR VGND sg13g2_mux2_1
X_2781_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[2\] net767 _0748_ _0528_
+ VPWR VGND sg13g2_mux2_1
X_4520_ _2143_ VPWR _2150_ VGND _0656_ _2139_ sg13g2_o21ai_1
X_4451_ tmds_green.n132 tmds_green.n126 net600 _2086_ VPWR VGND sg13g2_nand3_1
XFILLER_8_795 VPWR VGND sg13g2_fill_2
X_3402_ _1067_ _1068_ _1070_ _1071_ VPWR VGND sg13g2_or3_1
X_4382_ _2025_ _2024_ _2027_ VPWR VGND sg13g2_xor2_1
X_3333_ net745 _1021_ _0351_ VPWR VGND sg13g2_nor2_1
Xfanout708 net711 net708 VPWR VGND sg13g2_buf_8
Xfanout719 net723 net719 VPWR VGND sg13g2_buf_8
X_3264_ _0809_ _0966_ _0329_ VPWR VGND sg13g2_nor2_1
X_5003_ net237 VGND VPWR _0431_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[2\]
+ _0088_ sg13g2_dfrbpq_1
XFILLER_39_666 VPWR VGND sg13g2_decap_4
X_3195_ VGND VPWR _0917_ _0919_ _0278_ _0920_ sg13g2_a21oi_1
XFILLER_34_371 VPWR VGND sg13g2_fill_2
X_2979_ net775 _0796_ _0798_ VPWR VGND sg13g2_nor2_1
X_4718_ net667 net720 _0148_ VPWR VGND sg13g2_nor2_1
X_4649_ net669 net722 _0079_ VPWR VGND sg13g2_nor2_1
XFILLER_39_12 VPWR VGND sg13g2_decap_4
XFILLER_39_34 VPWR VGND sg13g2_decap_4
X_4900__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_29_121 VPWR VGND sg13g2_decap_4
XFILLER_45_603 VPWR VGND sg13g2_decap_8
XFILLER_33_809 VPWR VGND sg13g2_fill_2
XFILLER_38_1000 VPWR VGND sg13g2_decap_8
XFILLER_13_544 VPWR VGND sg13g2_fill_1
XFILLER_41_864 VPWR VGND sg13g2_fill_1
XFILLER_9_504 VPWR VGND sg13g2_decap_8
X_5152__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_40_396 VPWR VGND sg13g2_fill_2
XFILLER_49_931 VPWR VGND sg13g2_decap_8
X_3951_ _1619_ net613 _1618_ VPWR VGND sg13g2_nand2b_1
XFILLER_35_179 VPWR VGND sg13g2_fill_2
X_2902_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\] net755 _0778_ _0428_
+ VPWR VGND sg13g2_mux2_1
X_3882_ _1550_ VPWR _1551_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[2\]\[3\]
+ net553 sg13g2_o21ai_1
X_2833_ net762 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[2\] _0760_ _0479_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_363 VPWR VGND sg13g2_fill_1
X_2764_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[1\] _0742_ _0539_
+ VPWR VGND sg13g2_mux2_1
X_5014__216 VPWR VGND net216 sg13g2_tiehi
X_4503_ _2134_ tmds_blue.n132 _2133_ VPWR VGND sg13g2_xnor2_1
X_2695_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[0\] net793 _0724_ _0590_
+ VPWR VGND sg13g2_mux2_1
X_4434_ _2073_ net604 tmds_blue.n132 VPWR VGND sg13g2_xnor2_1
X_4365_ _0869_ tmds_red.dc_balancing_reg\[1\] _2001_ _2011_ VPWR VGND sg13g2_a21o_1
X_3316_ _1003_ VPWR _1006_ VGND _1004_ _1005_ sg13g2_o21ai_1
Xfanout549 _0682_ net549 VPWR VGND sg13g2_buf_8
X_4296_ VGND VPWR _1942_ _1956_ _1958_ _1925_ sg13g2_a21oi_1
X_3247_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[2\] videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\]
+ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[0\] _0955_ VPWR VGND sg13g2_or3_1
X_3178_ _0907_ _0903_ _0905_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_820 VPWR VGND sg13g2_decap_8
XFILLER_41_149 VPWR VGND sg13g2_fill_2
XFILLER_1_223 VPWR VGND sg13g2_fill_2
XFILLER_2_768 VPWR VGND sg13g2_decap_8
XFILLER_49_227 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_46_923 VPWR VGND sg13g2_decap_8
XFILLER_18_614 VPWR VGND sg13g2_fill_1
X_4861__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_17_124 VPWR VGND sg13g2_fill_2
XFILLER_18_647 VPWR VGND sg13g2_decap_4
XFILLER_18_658 VPWR VGND sg13g2_fill_2
XFILLER_18_669 VPWR VGND sg13g2_decap_8
XFILLER_33_606 VPWR VGND sg13g2_decap_8
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
X_4150_ _1807_ _1811_ _1812_ VPWR VGND sg13g2_nor2_1
X_3101_ green_tmds_par\[9\] net697 serialize.n428\[9\] VPWR VGND sg13g2_and2_1
X_4081_ _1746_ _1704_ _1739_ VPWR VGND sg13g2_nand2_1
X_3032_ _0807_ VPWR _0827_ VGND videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ _0822_ sg13g2_o21ai_1
X_4983_ net280 VGND VPWR _0411_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[2\]
+ _0068_ sg13g2_dfrbpq_1
XFILLER_20_801 VPWR VGND sg13g2_decap_4
X_3934_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\] net581 _1602_ VPWR
+ VGND sg13g2_nor2_1
X_3865_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\] net567 _1534_ VPWR
+ VGND sg13g2_nor2_1
X_2816_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[2\] net765 _0755_ _0491_
+ VPWR VGND sg13g2_mux2_1
X_3796_ _1465_ _0701_ _0650_ net593 _0635_ VPWR VGND sg13g2_a22oi_1
X_2747_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\] net759 _0739_ _0553_
+ VPWR VGND sg13g2_mux2_1
X_2678_ _0719_ _0718_ VPWR VGND net545 sg13g2_nand2b_2
X_4417_ _2058_ _2059_ _2060_ VPWR VGND sg13g2_and2_1
X_4348_ _1995_ tmds_red.n132 tmds_red.dc_balancing_reg\[1\] VPWR VGND sg13g2_xnor2_1
X_4279_ VPWR _1941_ _1940_ VGND sg13g2_inv_1
XFILLER_39_260 VPWR VGND sg13g2_fill_2
XFILLER_27_400 VPWR VGND sg13g2_decap_4
X_4882__85 VPWR VGND net85 sg13g2_tiehi
XFILLER_15_617 VPWR VGND sg13g2_fill_1
XFILLER_28_978 VPWR VGND sg13g2_decap_8
XFILLER_43_948 VPWR VGND sg13g2_decap_8
XFILLER_42_425 VPWR VGND sg13g2_fill_1
XFILLER_11_834 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_10_366 VPWR VGND sg13g2_decap_8
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_6_337 VPWR VGND sg13g2_fill_1
XFILLER_19_923 VPWR VGND sg13g2_decap_8
XFILLER_33_403 VPWR VGND sg13g2_decap_4
XFILLER_34_915 VPWR VGND sg13g2_decap_8
XFILLER_33_436 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_decap_8
X_3650_ videogen.test_lut_thingy.pixel_feeder_inst.row\[29\]\[2\] net568 _1319_ VPWR
+ VGND sg13g2_nor2_1
X_3581_ _1248_ _1249_ _1250_ VPWR VGND sg13g2_nor2_2
X_2601_ VPWR _0657_ tmds_blue.dc_balancing_reg\[3\] VGND sg13g2_inv_1
XFILLER_6_893 VPWR VGND sg13g2_decap_8
X_4202_ _1864_ _1846_ _1863_ VPWR VGND sg13g2_xnor2_1
X_5182_ net293 VGND VPWR _0606_ videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[0\]
+ _0254_ sg13g2_dfrbpq_1
XFILLER_3_72 VPWR VGND sg13g2_fill_2
X_4133_ _1398_ _1591_ _1700_ _1796_ VPWR VGND sg13g2_or3_1
X_4064_ _1729_ net544 _1708_ VPWR VGND sg13g2_xnor2_1
X_3015_ videogen.fancy_shader.video_x\[2\] _0810_ _0811_ VPWR VGND sg13g2_and2_1
XFILLER_37_775 VPWR VGND sg13g2_decap_8
XFILLER_37_753 VPWR VGND sg13g2_decap_4
X_4966_ net313 VGND VPWR _0394_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\]
+ _0051_ sg13g2_dfrbpq_1
X_4897_ net56 VGND VPWR _0325_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\]
+ net631 sg13g2_dfrbpq_2
XFILLER_20_620 VPWR VGND sg13g2_decap_8
X_3917_ net619 _1582_ _1584_ _1585_ _1586_ VPWR VGND sg13g2_nor4_1
X_3848_ net621 VPWR _1517_ VGND _1513_ _1516_ sg13g2_o21ai_1
X_3779_ net622 VPWR _1448_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\]
+ net587 sg13g2_o21ai_1
X_5066__264 VPWR VGND net264 sg13g2_tiehi
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_42_255 VPWR VGND sg13g2_fill_2
XFILLER_42_222 VPWR VGND sg13g2_decap_8
X_4870__99 VPWR VGND net99 sg13g2_tiehi
XFILLER_31_907 VPWR VGND sg13g2_decap_8
XFILLER_43_789 VPWR VGND sg13g2_decap_4
XFILLER_23_491 VPWR VGND sg13g2_fill_2
XFILLER_10_141 VPWR VGND sg13g2_decap_8
XFILLER_7_635 VPWR VGND sg13g2_fill_1
XFILLER_7_668 VPWR VGND sg13g2_fill_2
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_18_252 VPWR VGND sg13g2_fill_1
XFILLER_46_594 VPWR VGND sg13g2_decap_8
XFILLER_34_712 VPWR VGND sg13g2_decap_4
X_4820_ net652 net704 _0250_ VPWR VGND sg13g2_nor2_1
XFILLER_22_918 VPWR VGND sg13g2_decap_8
XFILLER_33_288 VPWR VGND sg13g2_fill_1
X_4751_ net673 net725 _0181_ VPWR VGND sg13g2_nor2_1
X_4682_ net675 net727 _0112_ VPWR VGND sg13g2_nor2_1
XFILLER_30_973 VPWR VGND sg13g2_decap_8
X_3702_ net612 VPWR _1371_ VGND _1365_ _1370_ sg13g2_o21ai_1
X_3633_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\] net585 _1302_ VPWR
+ VGND sg13g2_nor2_1
X_3564_ VGND VPWR _1233_ videogen.fancy_shader.video_x\[0\] net608 sg13g2_or2_1
X_3495_ _1164_ _1161_ _1162_ _1159_ _1127_ VPWR VGND sg13g2_a22oi_1
X_5234_ net799 VGND VPWR serialize.n429\[8\] serialize.n417\[6\] clknet_3_0__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4989__269 VPWR VGND net269 sg13g2_tiehi
X_5165_ net207 VGND VPWR _0589_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[3\]
+ _0237_ sg13g2_dfrbpq_1
X_4116_ _1754_ _1768_ _1779_ _1781_ VPWR VGND sg13g2_or3_1
X_5096_ net306 VGND VPWR _0520_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[2\]
+ _0168_ sg13g2_dfrbpq_1
X_4047_ _1710_ VPWR _1712_ VGND _1164_ _1165_ sg13g2_o21ai_1
XFILLER_24_222 VPWR VGND sg13g2_decap_8
X_4949_ net335 VGND VPWR _0377_ tmds_green.n126 net643 sg13g2_dfrbpq_2
XFILLER_33_47 VPWR VGND sg13g2_decap_4
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
XFILLER_20_472 VPWR VGND sg13g2_decap_4
XFILLER_3_159 VPWR VGND sg13g2_decap_8
X_4968__309 VPWR VGND net309 sg13g2_tiehi
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_837 VPWR VGND sg13g2_decap_8
XFILLER_47_314 VPWR VGND sg13g2_decap_4
XFILLER_43_575 VPWR VGND sg13g2_decap_8
XFILLER_16_778 VPWR VGND sg13g2_decap_8
XFILLER_12_940 VPWR VGND sg13g2_decap_8
XFILLER_15_299 VPWR VGND sg13g2_decap_8
XFILLER_30_225 VPWR VGND sg13g2_fill_1
XFILLER_30_247 VPWR VGND sg13g2_decap_4
XFILLER_8_933 VPWR VGND sg13g2_decap_8
X_3280_ videogen.test_lut_thingy.pixel_feeder_inst.h_counter\[1\] _0818_ _0977_ VPWR
+ VGND sg13g2_and2_1
XFILLER_39_804 VPWR VGND sg13g2_decap_4
XFILLER_24_4 VPWR VGND sg13g2_fill_1
XFILLER_47_892 VPWR VGND sg13g2_decap_8
XFILLER_34_520 VPWR VGND sg13g2_decap_8
XFILLER_34_564 VPWR VGND sg13g2_fill_2
X_4803_ net690 net741 _0233_ VPWR VGND sg13g2_nor2_1
X_4734_ net677 net729 _0164_ VPWR VGND sg13g2_nor2_1
X_2995_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[1\] net774 _0801_ _0284_
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_258 VPWR VGND sg13g2_decap_8
XFILLER_21_269 VPWR VGND sg13g2_decap_8
X_4665_ net685 net737 _0095_ VPWR VGND sg13g2_nor2_1
X_4596_ net665 net717 _0026_ VPWR VGND sg13g2_nor2_1
X_3616_ _1064_ _1281_ _1285_ VPWR VGND sg13g2_and2_1
X_3547_ _1216_ _1198_ _1200_ VPWR VGND sg13g2_nand2_1
X_3478_ _1147_ _1142_ _1145_ VPWR VGND sg13g2_xnor2_1
X_5217_ net804 VGND VPWR serialize.n428\[9\] serialize.n414\[7\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5148_ net385 VGND VPWR _0572_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[2\]
+ _0220_ sg13g2_dfrbpq_1
XFILLER_29_325 VPWR VGND sg13g2_decap_8
XFILLER_29_336 VPWR VGND sg13g2_fill_1
X_5079_ net379 VGND VPWR _0503_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[2\]
+ _0160_ sg13g2_dfrbpq_1
XFILLER_38_881 VPWR VGND sg13g2_decap_8
X_5104__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_13_704 VPWR VGND sg13g2_decap_4
XFILLER_9_708 VPWR VGND sg13g2_fill_2
XFILLER_12_236 VPWR VGND sg13g2_decap_8
XFILLER_9_719 VPWR VGND sg13g2_fill_2
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_0_641 VPWR VGND sg13g2_decap_8
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_48_634 VPWR VGND sg13g2_decap_4
XFILLER_44_851 VPWR VGND sg13g2_decap_8
XFILLER_44_862 VPWR VGND sg13g2_fill_1
X_2780_ videogen.test_lut_thingy.pixel_feeder_inst.row\[34\]\[3\] net757 _0748_ _0529_
+ VPWR VGND sg13g2_mux2_1
X_4450_ _2085_ net599 tmds_green.n126 VPWR VGND sg13g2_nand2_1
X_3401_ _1070_ videogen.fancy_shader.video_y\[4\] videogen.fancy_shader.n646\[4\]
+ VPWR VGND sg13g2_xnor2_1
X_4381_ _2024_ _2025_ _2026_ VPWR VGND sg13g2_and2_1
X_3332_ _1021_ videogen.fancy_shader.n646\[5\] _1019_ VPWR VGND sg13g2_xnor2_1
Xfanout709 net711 net709 VPWR VGND sg13g2_buf_8
X_3263_ _0965_ net610 _0966_ VPWR VGND sg13g2_xor2_1
XFILLER_39_645 VPWR VGND sg13g2_decap_8
X_5002_ net239 VGND VPWR _0430_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[1\]
+ _0087_ sg13g2_dfrbpq_1
XFILLER_22_1016 VPWR VGND sg13g2_decap_8
X_3194_ _0852_ VPWR _0920_ VGND _0917_ _0919_ sg13g2_o21ai_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
XFILLER_27_807 VPWR VGND sg13g2_fill_2
XFILLER_19_380 VPWR VGND sg13g2_decap_4
XFILLER_35_873 VPWR VGND sg13g2_decap_8
XFILLER_22_512 VPWR VGND sg13g2_decap_8
XFILLER_14_49 VPWR VGND sg13g2_decap_8
X_2978_ net764 videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\] _0796_ _0297_
+ VPWR VGND sg13g2_mux2_1
X_4717_ net660 net712 _0147_ VPWR VGND sg13g2_nor2_1
X_4648_ net669 net722 _0078_ VPWR VGND sg13g2_nor2_1
X_4579_ VGND VPWR _0882_ _0917_ _0277_ _0918_ sg13g2_a21oi_1
XFILLER_39_57 VPWR VGND sg13g2_fill_1
XFILLER_45_615 VPWR VGND sg13g2_fill_2
XFILLER_41_821 VPWR VGND sg13g2_fill_2
XFILLER_40_320 VPWR VGND sg13g2_decap_8
XFILLER_13_512 VPWR VGND sg13g2_decap_8
XFILLER_26_895 VPWR VGND sg13g2_decap_8
X_4978__290 VPWR VGND net290 sg13g2_tiehi
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_0_460 VPWR VGND sg13g2_decap_8
XFILLER_49_987 VPWR VGND sg13g2_decap_8
XFILLER_36_637 VPWR VGND sg13g2_decap_8
XFILLER_17_840 VPWR VGND sg13g2_fill_1
XFILLER_35_147 VPWR VGND sg13g2_fill_1
X_3950_ net597 _1612_ _1617_ _1618_ VPWR VGND sg13g2_nor3_1
X_2901_ _0728_ _0772_ _0778_ VPWR VGND sg13g2_nor2_2
XFILLER_32_843 VPWR VGND sg13g2_decap_8
X_3881_ _1550_ _0701_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_31_342 VPWR VGND sg13g2_fill_2
X_2832_ net753 videogen.test_lut_thingy.pixel_feeder_inst.row\[8\]\[3\] _0760_ _0480_
+ VPWR VGND sg13g2_mux2_1
X_2763_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[2\] _0742_ _0540_
+ VPWR VGND sg13g2_mux2_1
X_4502_ _2133_ tmds_blue.n193 tmds_blue.dc_balancing_reg\[1\] VPWR VGND sg13g2_xnor2_1
XFILLER_8_593 VPWR VGND sg13g2_decap_8
X_2694_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[1\] net782 _0724_ _0591_
+ VPWR VGND sg13g2_mux2_1
X_4433_ VGND VPWR net605 _2072_ _0615_ _2069_ sg13g2_a21oi_1
X_4364_ VGND VPWR _2007_ _2009_ _2010_ _0911_ sg13g2_a21oi_1
X_3315_ _1005_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_x\[1\]
+ VPWR VGND sg13g2_xnor2_1
X_4295_ _1957_ _1925_ _1942_ _1956_ VPWR VGND sg13g2_and3_1
X_3246_ VPWR _0323_ _0954_ VGND sg13g2_inv_1
XFILLER_39_431 VPWR VGND sg13g2_decap_4
X_3177_ _0906_ _0903_ _0905_ _0866_ _0664_ VPWR VGND sg13g2_a22oi_1
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_41_36 VPWR VGND sg13g2_fill_2
XFILLER_6_508 VPWR VGND sg13g2_decap_4
XFILLER_22_397 VPWR VGND sg13g2_fill_1
XFILLER_49_206 VPWR VGND sg13g2_decap_8
XFILLER_46_902 VPWR VGND sg13g2_decap_8
XFILLER_46_979 VPWR VGND sg13g2_decap_8
XFILLER_14_810 VPWR VGND sg13g2_fill_2
XFILLER_14_832 VPWR VGND sg13g2_fill_2
XFILLER_41_662 VPWR VGND sg13g2_fill_2
XFILLER_9_324 VPWR VGND sg13g2_decap_8
XFILLER_40_183 VPWR VGND sg13g2_decap_8
XFILLER_5_541 VPWR VGND sg13g2_fill_2
XFILLER_31_91 VPWR VGND sg13g2_fill_1
XFILLER_5_585 VPWR VGND sg13g2_fill_1
X_3100_ green_tmds_par\[8\] net695 serialize.n428\[8\] VPWR VGND sg13g2_and2_1
X_4080_ _1745_ _1707_ _1742_ VPWR VGND sg13g2_xnor2_1
X_3031_ VGND VPWR _0808_ _0826_ _0002_ _0371_ sg13g2_a21oi_1
XFILLER_36_401 VPWR VGND sg13g2_decap_8
XFILLER_36_412 VPWR VGND sg13g2_fill_1
XFILLER_36_434 VPWR VGND sg13g2_decap_8
XFILLER_37_979 VPWR VGND sg13g2_decap_8
X_4982_ net282 VGND VPWR _0410_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\]
+ _0067_ sg13g2_dfrbpq_1
X_3933_ _1597_ _1598_ _1599_ _1600_ _1601_ VPWR VGND sg13g2_nor4_1
XFILLER_16_191 VPWR VGND sg13g2_fill_2
X_3864_ _1532_ VPWR _1533_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[41\]\[3\]
+ net566 sg13g2_o21ai_1
X_5199__65 VPWR VGND net65 sg13g2_tiehi
X_2815_ videogen.test_lut_thingy.pixel_feeder_inst.row\[3\]\[3\] net754 _0755_ _0492_
+ VPWR VGND sg13g2_mux2_1
X_3795_ net621 VPWR _1464_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[1\]
+ net563 sg13g2_o21ai_1
X_2746_ _0726_ _0733_ _0739_ VPWR VGND sg13g2_nor2_2
X_2677_ _0693_ _0696_ _0718_ VPWR VGND sg13g2_nor2_2
X_4416_ _0655_ _2056_ tmds_blue.n193 _2059_ VPWR VGND sg13g2_nand3_1
X_4347_ tmds_red.dc_balancing_reg\[0\] _0852_ _0509_ VPWR VGND sg13g2_and2_1
X_5168__183 VPWR VGND net183 sg13g2_tiehi
X_4278_ VGND VPWR _1940_ _1939_ _1922_ sg13g2_or2_1
X_3229_ _0943_ net796 _0942_ VPWR VGND sg13g2_nand2_2
XFILLER_28_957 VPWR VGND sg13g2_decap_8
XFILLER_43_905 VPWR VGND sg13g2_fill_1
XFILLER_36_69 VPWR VGND sg13g2_decap_4
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_23_640 VPWR VGND sg13g2_decap_8
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_11_813 VPWR VGND sg13g2_fill_2
XFILLER_7_806 VPWR VGND sg13g2_decap_4
XFILLER_6_327 VPWR VGND sg13g2_fill_2
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_46_743 VPWR VGND sg13g2_decap_8
XFILLER_18_467 VPWR VGND sg13g2_fill_1
XFILLER_18_478 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_9_132 VPWR VGND sg13g2_decap_4
X_3580_ _1146_ _1246_ _1249_ VPWR VGND sg13g2_nor2_1
X_2600_ VPWR _0656_ tmds_blue.dc_balancing_reg\[1\] VGND sg13g2_inv_1
XFILLER_6_872 VPWR VGND sg13g2_decap_8
XFILLER_6_850 VPWR VGND sg13g2_fill_2
X_4201_ _1849_ VPWR _1863_ VGND _1853_ _1855_ sg13g2_o21ai_1
X_5181_ net308 VGND VPWR _0605_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\]
+ _0253_ sg13g2_dfrbpq_1
X_4132_ _1795_ _1496_ _1591_ VPWR VGND sg13g2_nand2_1
X_4063_ _1725_ _1727_ _1728_ VPWR VGND sg13g2_and2_1
X_3014_ videogen.fancy_shader.video_x\[1\] videogen.fancy_shader.video_x\[0\] _0810_
+ VPWR VGND sg13g2_and2_1
XFILLER_36_253 VPWR VGND sg13g2_decap_8
XFILLER_25_949 VPWR VGND sg13g2_decap_8
X_4965_ net315 VGND VPWR _0393_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[0\]
+ _0050_ sg13g2_dfrbpq_1
X_3916_ videogen.test_lut_thingy.pixel_feeder_inst.row\[25\]\[3\] net565 _1585_ VPWR
+ VGND sg13g2_nor2_1
X_4896_ net58 VGND VPWR _0324_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[0\]
+ net630 sg13g2_dfrbpq_2
X_3847_ _1515_ VPWR _1516_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[60\]\[3\]
+ net586 sg13g2_o21ai_1
X_3778_ _1446_ VPWR _1447_ VGND _1410_ _1422_ sg13g2_o21ai_1
X_2729_ net788 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[0\] _0734_ _0566_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_426 VPWR VGND sg13g2_fill_2
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_27_275 VPWR VGND sg13g2_fill_1
XFILLER_43_746 VPWR VGND sg13g2_fill_1
XFILLER_42_234 VPWR VGND sg13g2_decap_8
XFILLER_11_665 VPWR VGND sg13g2_fill_1
XFILLER_6_135 VPWR VGND sg13g2_fill_2
X_5114__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_3_864 VPWR VGND sg13g2_decap_8
XFILLER_2_352 VPWR VGND sg13g2_decap_8
X_4914__394 VPWR VGND net394 sg13g2_tiehi
X_5084__365 VPWR VGND net365 sg13g2_tiehi
XFILLER_19_776 VPWR VGND sg13g2_fill_2
XFILLER_18_264 VPWR VGND sg13g2_decap_4
XFILLER_33_245 VPWR VGND sg13g2_decap_4
XFILLER_15_982 VPWR VGND sg13g2_decap_8
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
X_4750_ net673 net725 _0180_ VPWR VGND sg13g2_nor2_1
X_4681_ net676 net728 _0111_ VPWR VGND sg13g2_nor2_1
XFILLER_30_952 VPWR VGND sg13g2_decap_8
X_3701_ net622 VPWR _1370_ VGND _1366_ _1369_ sg13g2_o21ai_1
X_3632_ net614 VPWR _1301_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[2\]
+ net552 sg13g2_o21ai_1
X_3563_ _1232_ _1063_ _1231_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_3494_ _1163_ _1161_ _1162_ VPWR VGND sg13g2_nand2_1
X_5233_ net799 VGND VPWR serialize.n429\[7\] serialize.n417\[5\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5164_ net215 VGND VPWR _0588_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[2\]
+ _0236_ sg13g2_dfrbpq_1
X_4115_ _1754_ VPWR _1780_ VGND _1768_ _1779_ sg13g2_o21ai_1
XFILLER_29_507 VPWR VGND sg13g2_decap_8
X_5095_ net310 VGND VPWR _0519_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[1\]
+ _0167_ sg13g2_dfrbpq_1
X_4046_ _1164_ _1165_ _1710_ _1711_ VPWR VGND sg13g2_or3_1
XFILLER_37_573 VPWR VGND sg13g2_decap_4
XFILLER_25_702 VPWR VGND sg13g2_fill_1
XFILLER_13_919 VPWR VGND sg13g2_decap_8
XFILLER_12_429 VPWR VGND sg13g2_decap_8
X_4948_ net336 VGND VPWR _0376_ tmds_green.n100 net636 sg13g2_dfrbpq_2
XFILLER_33_790 VPWR VGND sg13g2_decap_4
X_4879_ net89 VGND VPWR _0307_ videogen.fancy_shader.video_x\[8\] net634 sg13g2_dfrbpq_2
XFILLER_20_451 VPWR VGND sg13g2_fill_2
XFILLER_21_985 VPWR VGND sg13g2_decap_8
XFILLER_4_628 VPWR VGND sg13g2_decap_8
XFILLER_0_845 VPWR VGND sg13g2_decap_8
XFILLER_48_816 VPWR VGND sg13g2_decap_8
XFILLER_28_573 VPWR VGND sg13g2_decap_8
XFILLER_15_223 VPWR VGND sg13g2_decap_4
XFILLER_15_234 VPWR VGND sg13g2_fill_2
XFILLER_16_746 VPWR VGND sg13g2_fill_1
XFILLER_15_267 VPWR VGND sg13g2_decap_8
XFILLER_8_912 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_8_989 VPWR VGND sg13g2_decap_8
XFILLER_7_477 VPWR VGND sg13g2_decap_8
X_4988__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_39_849 VPWR VGND sg13g2_fill_1
XFILLER_39_838 VPWR VGND sg13g2_decap_8
X_5045__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_17_4 VPWR VGND sg13g2_decap_8
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_41 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_74 VPWR VGND sg13g2_fill_1
X_4841__149 VPWR VGND net149 sg13g2_tiehi
X_4802_ net691 net741 _0232_ VPWR VGND sg13g2_nor2_1
X_2994_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[2\] net763 _0801_ _0285_
+ VPWR VGND sg13g2_mux2_1
X_4733_ net677 net729 _0163_ VPWR VGND sg13g2_nor2_1
X_4664_ net684 net736 _0094_ VPWR VGND sg13g2_nor2_1
X_4595_ net649 net703 _0025_ VPWR VGND sg13g2_nor2_1
X_3615_ VGND VPWR _1281_ _1283_ _1284_ _1064_ sg13g2_a21oi_1
X_3546_ _1212_ _1214_ _1208_ _1215_ VPWR VGND sg13g2_nand3_1
X_5216_ net801 VGND VPWR serialize.n428\[8\] serialize.n414\[6\] clknet_3_1__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_3477_ _1145_ _1142_ _1146_ VPWR VGND sg13g2_xor2_1
X_5147_ net393 VGND VPWR _0571_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[1\]
+ _0219_ sg13g2_dfrbpq_1
XFILLER_28_48 VPWR VGND sg13g2_fill_1
X_5078_ net383 VGND VPWR _0502_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[1\]
+ _0159_ sg13g2_dfrbpq_1
XFILLER_28_59 VPWR VGND sg13g2_fill_1
XFILLER_38_860 VPWR VGND sg13g2_fill_2
X_4029_ VGND VPWR _1299_ _1696_ _0374_ _1596_ sg13g2_a21oi_1
XFILLER_37_381 VPWR VGND sg13g2_fill_2
XFILLER_12_215 VPWR VGND sg13g2_decap_8
XFILLER_40_546 VPWR VGND sg13g2_decap_4
XFILLER_21_793 VPWR VGND sg13g2_decap_4
XFILLER_5_937 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_30 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_35_329 VPWR VGND sg13g2_fill_2
XFILLER_43_384 VPWR VGND sg13g2_fill_1
XFILLER_34_91 VPWR VGND sg13g2_fill_2
XFILLER_15_1024 VPWR VGND sg13g2_decap_4
XFILLER_8_764 VPWR VGND sg13g2_decap_4
XFILLER_11_270 VPWR VGND sg13g2_fill_2
XFILLER_11_281 VPWR VGND sg13g2_decap_8
XFILLER_8_797 VPWR VGND sg13g2_fill_1
X_3400_ _1069_ videogen.fancy_shader.video_y\[4\] videogen.fancy_shader.n646\[4\]
+ VPWR VGND sg13g2_nand2_1
X_4380_ _2025_ _0907_ _1998_ VPWR VGND sg13g2_nand2_1
XFILLER_4_981 VPWR VGND sg13g2_decap_8
X_3331_ net750 _1019_ _1020_ _0350_ VPWR VGND sg13g2_nor3_1
X_3262_ _0328_ _0808_ _0964_ _0965_ VPWR VGND sg13g2_and3_1
X_5001_ net241 VGND VPWR _0429_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\]
+ _0086_ sg13g2_dfrbpq_1
X_3193_ _0919_ _0663_ _0875_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_852 VPWR VGND sg13g2_decap_4
XFILLER_35_885 VPWR VGND sg13g2_decap_4
XFILLER_14_17 VPWR VGND sg13g2_fill_2
XFILLER_34_373 VPWR VGND sg13g2_fill_1
XFILLER_34_395 VPWR VGND sg13g2_fill_2
XFILLER_14_28 VPWR VGND sg13g2_decap_8
X_2977_ VGND VPWR _0649_ _0796_ _0298_ _0797_ sg13g2_a21oi_1
X_4716_ net660 net712 _0146_ VPWR VGND sg13g2_nor2_1
X_4647_ net670 net721 _0077_ VPWR VGND sg13g2_nor2_1
XFILLER_30_16 VPWR VGND sg13g2_decap_4
XFILLER_30_49 VPWR VGND sg13g2_fill_2
X_4578_ _0654_ net571 _0272_ VPWR VGND sg13g2_nor2_1
XFILLER_2_929 VPWR VGND sg13g2_decap_8
X_3529_ _1188_ _1197_ _1187_ _1198_ VPWR VGND sg13g2_nand3_1
XFILLER_45_649 VPWR VGND sg13g2_fill_1
XFILLER_45_638 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_4
XFILLER_44_148 VPWR VGND sg13g2_fill_2
XFILLER_26_874 VPWR VGND sg13g2_decap_8
XFILLER_25_362 VPWR VGND sg13g2_decap_8
XFILLER_41_855 VPWR VGND sg13g2_decap_8
XFILLER_4_233 VPWR VGND sg13g2_fill_2
XFILLER_5_778 VPWR VGND sg13g2_fill_1
XFILLER_20_71 VPWR VGND sg13g2_decap_4
XFILLER_1_984 VPWR VGND sg13g2_decap_8
XFILLER_49_966 VPWR VGND sg13g2_decap_8
XFILLER_0_494 VPWR VGND sg13g2_decap_8
XFILLER_35_115 VPWR VGND sg13g2_decap_4
X_2900_ videogen.test_lut_thingy.pixel_feeder_inst.row\[52\]\[0\] net788 _0777_ _0429_
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_373 VPWR VGND sg13g2_decap_8
XFILLER_31_310 VPWR VGND sg13g2_decap_4
X_3880_ videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[3\] net586 _1549_ VPWR
+ VGND sg13g2_nor2_1
X_2831_ _0760_ _0699_ _0720_ VPWR VGND sg13g2_nand2_2
X_2762_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[31\]\[3\] _0742_ _0541_
+ VPWR VGND sg13g2_mux2_1
X_4501_ net751 clockdiv.q0 net406 _0623_ VPWR VGND sg13g2_nor3_1
X_4432_ _2071_ _2070_ _2072_ VPWR VGND sg13g2_xor2_1
X_2693_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[2\] net770 _0724_ _0592_
+ VPWR VGND sg13g2_mux2_1
X_4363_ _2008_ VPWR _2009_ VGND net548 _1996_ sg13g2_o21ai_1
X_3314_ _1004_ videogen.fancy_shader.n646\[0\] videogen.fancy_shader.video_x\[0\]
+ VPWR VGND sg13g2_nand2_1
X_4294_ _1943_ VPWR _1956_ VGND _1944_ _1954_ sg13g2_o21ai_1
X_4894__62 VPWR VGND net62 sg13g2_tiehi
X_3245_ _0953_ VPWR _0954_ VGND videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ _0952_ sg13g2_o21ai_1
XFILLER_27_616 VPWR VGND sg13g2_decap_8
X_3176_ _0869_ _0904_ _0905_ VPWR VGND sg13g2_and2_1
XFILLER_26_104 VPWR VGND sg13g2_decap_8
XFILLER_41_129 VPWR VGND sg13g2_fill_2
XFILLER_22_310 VPWR VGND sg13g2_fill_1
XFILLER_25_49 VPWR VGND sg13g2_fill_2
XFILLER_34_170 VPWR VGND sg13g2_decap_8
XFILLER_22_321 VPWR VGND sg13g2_fill_2
XFILLER_34_181 VPWR VGND sg13g2_fill_2
XFILLER_41_48 VPWR VGND sg13g2_decap_8
XFILLER_2_737 VPWR VGND sg13g2_decap_4
XFILLER_45_402 VPWR VGND sg13g2_fill_1
XFILLER_46_958 VPWR VGND sg13g2_decap_8
XFILLER_40_162 VPWR VGND sg13g2_decap_4
XFILLER_13_365 VPWR VGND sg13g2_decap_8
XFILLER_9_336 VPWR VGND sg13g2_fill_2
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_5_564 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_1_781 VPWR VGND sg13g2_decap_8
XFILLER_49_741 VPWR VGND sg13g2_fill_2
X_3030_ _0822_ _0823_ net795 _0826_ VPWR VGND _0824_ sg13g2_nand4_1
XFILLER_24_619 VPWR VGND sg13g2_decap_8
XFILLER_36_468 VPWR VGND sg13g2_decap_8
XFILLER_45_991 VPWR VGND sg13g2_decap_8
X_4981_ net284 VGND VPWR _0409_ videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[0\]
+ _0066_ sg13g2_dfrbpq_1
X_4924__374 VPWR VGND net374 sg13g2_tiehi
X_3932_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[0\] net569 _1600_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_16_170 VPWR VGND sg13g2_fill_1
X_3863_ _1529_ _1530_ _1531_ _1532_ VPWR VGND sg13g2_nor3_1
X_2814_ _0714_ _0737_ _0755_ VPWR VGND sg13g2_nor2_2
XFILLER_31_173 VPWR VGND sg13g2_decap_8
X_3794_ net621 _1459_ _1460_ _1462_ _1463_ VPWR VGND sg13g2_nor4_1
XFILLER_8_391 VPWR VGND sg13g2_fill_1
XFILLER_11_29 VPWR VGND sg13g2_fill_1
X_2745_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[0\] net785 _0738_ _0554_
+ VPWR VGND sg13g2_mux2_1
X_2676_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[0\] net784 _0717_ _0602_
+ VPWR VGND sg13g2_mux2_1
X_4415_ _2058_ tmds_blue.dc_balancing_reg\[4\] tmds_blue.n193 VPWR VGND sg13g2_nand2b_1
X_4346_ VGND VPWR _0859_ _1994_ _0508_ net748 sg13g2_a21oi_1
X_4277_ VGND VPWR _1912_ _1916_ _1939_ _1921_ sg13g2_a21oi_1
X_3228_ _0942_ _0677_ _0683_ VPWR VGND sg13g2_nand2_2
XFILLER_39_284 VPWR VGND sg13g2_decap_4
X_3159_ _0888_ tmds_red.n100 _0869_ VPWR VGND sg13g2_nand2_1
XFILLER_28_936 VPWR VGND sg13g2_decap_8
XFILLER_27_446 VPWR VGND sg13g2_fill_2
XFILLER_22_140 VPWR VGND sg13g2_decap_8
XFILLER_2_567 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_fill_2
XFILLER_18_413 VPWR VGND sg13g2_decap_8
XFILLER_19_958 VPWR VGND sg13g2_decap_8
XFILLER_27_991 VPWR VGND sg13g2_decap_8
XFILLER_14_674 VPWR VGND sg13g2_fill_2
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_fill_1
X_4200_ VGND VPWR _1862_ _1861_ _1853_ sg13g2_or2_1
X_5180_ net347 VGND VPWR _0604_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\]
+ _0252_ sg13g2_dfrbpq_1
XFILLER_3_74 VPWR VGND sg13g2_fill_1
X_4131_ _1792_ _1794_ _1790_ _0376_ VPWR VGND sg13g2_nand3_1
X_4062_ _1718_ VPWR _1727_ VGND _1721_ _1722_ sg13g2_o21ai_1
XFILLER_3_85 VPWR VGND sg13g2_fill_1
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
X_3013_ _0809_ net795 VPWR VGND videogen.test_lut_thingy.pixel_feeder_inst.state\[0\]
+ sg13g2_nand2b_2
XFILLER_24_405 VPWR VGND sg13g2_fill_2
XFILLER_25_928 VPWR VGND sg13g2_decap_8
XFILLER_36_265 VPWR VGND sg13g2_decap_4
XFILLER_36_287 VPWR VGND sg13g2_decap_8
X_4964_ net317 VGND VPWR _0392_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\]
+ _0049_ sg13g2_dfrbpq_1
XFILLER_24_449 VPWR VGND sg13g2_fill_2
X_3915_ _1583_ VPWR _1584_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\]
+ net585 sg13g2_o21ai_1
X_4895_ net60 VGND VPWR _0323_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\]
+ net631 sg13g2_dfrbpq_2
XFILLER_32_493 VPWR VGND sg13g2_decap_4
XFILLER_33_994 VPWR VGND sg13g2_decap_8
XFILLER_22_17 VPWR VGND sg13g2_fill_2
X_3846_ VGND VPWR _0649_ _0701_ _1515_ _1514_ sg13g2_a21oi_1
XFILLER_20_677 VPWR VGND sg13g2_fill_2
XFILLER_20_699 VPWR VGND sg13g2_decap_8
X_3777_ net610 _1445_ _1446_ VPWR VGND sg13g2_nor2_1
XFILLER_3_309 VPWR VGND sg13g2_fill_1
X_2728_ net777 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\] _0734_ _0567_
+ VPWR VGND sg13g2_mux2_1
X_2659_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[0\] net784 _0708_ _0628_
+ VPWR VGND sg13g2_mux2_1
X_4329_ net747 _1984_ _0385_ VPWR VGND sg13g2_nor2_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_700 VPWR VGND sg13g2_fill_1
XFILLER_47_58 VPWR VGND sg13g2_fill_1
XFILLER_16_917 VPWR VGND sg13g2_decap_8
XFILLER_28_755 VPWR VGND sg13g2_decap_8
XFILLER_43_725 VPWR VGND sg13g2_decap_8
XFILLER_43_703 VPWR VGND sg13g2_fill_2
XFILLER_15_438 VPWR VGND sg13g2_fill_1
XFILLER_24_983 VPWR VGND sg13g2_decap_8
XFILLER_30_408 VPWR VGND sg13g2_decap_8
XFILLER_11_699 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_fill_2
XFILLER_3_843 VPWR VGND sg13g2_decap_8
XFILLER_2_320 VPWR VGND sg13g2_fill_1
Xfanout690 net691 net690 VPWR VGND sg13g2_buf_8
XFILLER_19_711 VPWR VGND sg13g2_decap_4
XFILLER_19_744 VPWR VGND sg13g2_decap_8
X_5121__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_46_563 VPWR VGND sg13g2_decap_8
XFILLER_34_747 VPWR VGND sg13g2_decap_4
XFILLER_15_961 VPWR VGND sg13g2_decap_8
XFILLER_30_931 VPWR VGND sg13g2_decap_8
X_3700_ _1368_ VPWR _1369_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[63\]\[2\]
+ net575 sg13g2_o21ai_1
XFILLER_41_290 VPWR VGND sg13g2_fill_1
X_4680_ net676 net728 _0110_ VPWR VGND sg13g2_nor2_1
X_3631_ _1300_ videogen.test_lut_thingy.pixel_feeder_inst.h_pix\[1\] _0647_ VPWR VGND
+ sg13g2_nand2_2
X_3562_ _1227_ _1230_ _1231_ VPWR VGND sg13g2_and2_1
X_3493_ _1103_ _1101_ _1104_ _1162_ VPWR VGND sg13g2_a21o_2
X_5232_ net800 VGND VPWR serialize.n429\[6\] serialize.n417\[4\] clknet_3_0__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_5163_ net223 VGND VPWR _0587_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[1\]
+ _0235_ sg13g2_dfrbpq_1
X_4114_ _1703_ _1770_ _1777_ _1779_ VPWR VGND sg13g2_nor3_1
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
X_5094_ net314 VGND VPWR _0518_ videogen.test_lut_thingy.pixel_feeder_inst.row\[36\]\[0\]
+ _0166_ sg13g2_dfrbpq_1
XFILLER_49_390 VPWR VGND sg13g2_decap_8
X_4045_ _1100_ _1709_ _1710_ VPWR VGND sg13g2_and2_1
XFILLER_17_17 VPWR VGND sg13g2_decap_4
XFILLER_25_714 VPWR VGND sg13g2_decap_8
XFILLER_12_408 VPWR VGND sg13g2_fill_1
X_4947_ net337 VGND VPWR _0375_ tmds_blue.n132 net636 sg13g2_dfrbpq_2
X_4878_ net90 VGND VPWR _0306_ videogen.fancy_shader.video_x\[7\] net634 sg13g2_dfrbpq_1
XFILLER_21_964 VPWR VGND sg13g2_decap_8
X_3829_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\] net553 _1498_ VPWR
+ VGND sg13g2_nor2_1
X_4907__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_0_824 VPWR VGND sg13g2_decap_8
X_5148__385 VPWR VGND net385 sg13g2_tiehi
XFILLER_47_305 VPWR VGND sg13g2_decap_4
XFILLER_43_511 VPWR VGND sg13g2_fill_2
XFILLER_43_555 VPWR VGND sg13g2_decap_8
XFILLER_31_706 VPWR VGND sg13g2_fill_2
XFILLER_31_739 VPWR VGND sg13g2_decap_8
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_8_968 VPWR VGND sg13g2_decap_8
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_4
XFILLER_47_850 VPWR VGND sg13g2_decap_8
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_decap_8
XFILLER_22_706 VPWR VGND sg13g2_fill_2
XFILLER_34_566 VPWR VGND sg13g2_fill_1
X_4801_ net691 net741 _0231_ VPWR VGND sg13g2_nor2_1
X_2993_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\] net756 _0801_ _0286_
+ VPWR VGND sg13g2_mux2_1
X_4995__253 VPWR VGND net253 sg13g2_tiehi
X_4732_ net677 net729 _0162_ VPWR VGND sg13g2_nor2_1
X_4663_ net684 net736 _0093_ VPWR VGND sg13g2_nor2_1
XFILLER_30_761 VPWR VGND sg13g2_decap_4
X_3614_ _1283_ _1275_ _1282_ VPWR VGND sg13g2_nand2_1
X_4594_ net649 net701 _0024_ VPWR VGND sg13g2_nor2_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_3545_ _1065_ _1189_ _1214_ VPWR VGND sg13g2_nor2_1
X_3476_ _1143_ _1144_ _1145_ VPWR VGND sg13g2_and2_1
X_5215_ net803 VGND VPWR serialize.n428\[7\] serialize.n414\[5\] clknet_3_7__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_4967__311 VPWR VGND net311 sg13g2_tiehi
X_5146_ net401 VGND VPWR _0570_ videogen.test_lut_thingy.pixel_feeder_inst.row\[23\]\[0\]
+ _0218_ sg13g2_dfrbpq_1
XFILLER_28_27 VPWR VGND sg13g2_decap_8
X_5077_ net387 VGND VPWR _0501_ videogen.test_lut_thingy.pixel_feeder_inst.row\[13\]\[0\]
+ _0158_ sg13g2_dfrbpq_1
X_4028_ VPWR _1696_ _1695_ VGND sg13g2_inv_1
XFILLER_25_522 VPWR VGND sg13g2_fill_1
XFILLER_25_566 VPWR VGND sg13g2_decap_4
XFILLER_40_525 VPWR VGND sg13g2_decap_8
XFILLER_40_503 VPWR VGND sg13g2_fill_2
XFILLER_13_728 VPWR VGND sg13g2_fill_2
XFILLER_20_282 VPWR VGND sg13g2_decap_4
XFILLER_5_916 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_20 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_4_459 VPWR VGND sg13g2_fill_2
XFILLER_0_698 VPWR VGND sg13g2_decap_8
XFILLER_28_360 VPWR VGND sg13g2_decap_8
XFILLER_29_883 VPWR VGND sg13g2_decap_4
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_31_525 VPWR VGND sg13g2_fill_1
XFILLER_15_1003 VPWR VGND sg13g2_decap_8
XFILLER_8_732 VPWR VGND sg13g2_fill_2
XFILLER_8_721 VPWR VGND sg13g2_decap_4
XFILLER_8_743 VPWR VGND sg13g2_decap_4
XFILLER_12_794 VPWR VGND sg13g2_fill_2
XFILLER_4_960 VPWR VGND sg13g2_decap_8
X_3330_ VGND VPWR videogen.fancy_shader.n646\[3\] _0996_ _1020_ videogen.fancy_shader.n646\[4\]
+ sg13g2_a21oi_1
X_5000_ net243 VGND VPWR _0428_ videogen.test_lut_thingy.pixel_feeder_inst.row\[53\]\[3\]
+ _0085_ sg13g2_dfrbpq_1
XFILLER_3_492 VPWR VGND sg13g2_decap_4
X_3261_ _0965_ net611 _0963_ VPWR VGND sg13g2_nand2_1
X_3192_ VGND VPWR _0882_ _0917_ _0276_ _0918_ sg13g2_a21oi_1
XFILLER_38_124 VPWR VGND sg13g2_decap_4
XFILLER_22_569 VPWR VGND sg13g2_decap_4
X_2976_ net754 _0796_ _0797_ VPWR VGND sg13g2_nor2_1
X_4715_ net678 net729 _0145_ VPWR VGND sg13g2_nor2_1
XFILLER_30_580 VPWR VGND sg13g2_decap_8
X_4646_ net670 net721 _0076_ VPWR VGND sg13g2_nor2_1
X_4577_ net677 net729 _0009_ VPWR VGND sg13g2_nor2_1
X_4934__354 VPWR VGND net354 sg13g2_tiehi
XFILLER_2_908 VPWR VGND sg13g2_decap_8
X_3528_ _1178_ _1195_ _1197_ VPWR VGND sg13g2_nor2_1
XFILLER_39_48 VPWR VGND sg13g2_decap_8
X_3459_ videogen.fancy_shader.video_x\[9\] videogen.fancy_shader.n646\[9\] _1128_
+ VPWR VGND sg13g2_xor2_1
X_5129_ net173 VGND VPWR _0553_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[3\]
+ _0201_ sg13g2_dfrbpq_1
XFILLER_45_617 VPWR VGND sg13g2_fill_1
XFILLER_38_1014 VPWR VGND sg13g2_decap_8
XFILLER_25_330 VPWR VGND sg13g2_fill_2
XFILLER_25_352 VPWR VGND sg13g2_fill_2
XFILLER_26_853 VPWR VGND sg13g2_decap_8
XFILLER_41_834 VPWR VGND sg13g2_decap_8
XFILLER_41_823 VPWR VGND sg13g2_fill_1
XFILLER_25_396 VPWR VGND sg13g2_decap_8
XFILLER_5_713 VPWR VGND sg13g2_fill_2
XFILLER_5_757 VPWR VGND sg13g2_fill_2
XFILLER_5_746 VPWR VGND sg13g2_fill_2
XFILLER_4_201 VPWR VGND sg13g2_decap_8
XFILLER_1_963 VPWR VGND sg13g2_decap_8
XFILLER_49_945 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_fill_1
XFILLER_36_606 VPWR VGND sg13g2_decap_8
XFILLER_32_812 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_fill_2
X_2830_ net789 videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[0\] _0759_ _0481_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_333 VPWR VGND sg13g2_decap_4
XFILLER_31_344 VPWR VGND sg13g2_fill_1
X_2761_ _0742_ _0716_ _0732_ VPWR VGND sg13g2_nand2_2
XFILLER_31_399 VPWR VGND sg13g2_fill_2
X_4500_ net572 _2132_ _0622_ VPWR VGND sg13g2_nor2_1
X_2692_ videogen.test_lut_thingy.pixel_feeder_inst.row\[18\]\[3\] net760 _0724_ _0593_
+ VPWR VGND sg13g2_mux2_1
X_4431_ _2071_ tmds_blue.n126 _2066_ VPWR VGND sg13g2_xnor2_1
X_4362_ _2004_ _1996_ _2008_ VPWR VGND sg13g2_xor2_1
X_3313_ _1003_ videogen.fancy_shader.n646\[1\] videogen.fancy_shader.video_x\[1\]
+ VPWR VGND sg13g2_nand2_1
X_4293_ VGND VPWR _1955_ _1954_ _1944_ sg13g2_or2_1
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
X_3244_ VGND VPWR videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[5\] _0952_ _0953_
+ _0943_ sg13g2_a21oi_1
XFILLER_6_1023 VPWR VGND sg13g2_fill_2
X_3175_ _0898_ _0888_ _0904_ VPWR VGND sg13g2_xor2_1
XFILLER_22_333 VPWR VGND sg13g2_fill_1
X_2959_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[0\] net793 _0792_ _0342_
+ VPWR VGND sg13g2_mux2_1
X_4629_ net652 net704 _0059_ VPWR VGND sg13g2_nor2_1
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_46_937 VPWR VGND sg13g2_decap_8
XFILLER_14_812 VPWR VGND sg13g2_fill_1
XFILLER_14_834 VPWR VGND sg13g2_fill_1
XFILLER_25_171 VPWR VGND sg13g2_fill_1
XFILLER_40_152 VPWR VGND sg13g2_decap_4
XFILLER_13_355 VPWR VGND sg13g2_fill_2
X_5156__281 VPWR VGND net281 sg13g2_tiehi
X_5117__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
X_5187__219 VPWR VGND net219 sg13g2_tiehi
XFILLER_5_543 VPWR VGND sg13g2_fill_1
Xoutput3 net3 tmds_b VPWR VGND sg13g2_buf_1
XFILLER_1_760 VPWR VGND sg13g2_decap_8
XFILLER_37_904 VPWR VGND sg13g2_fill_2
X_4980_ net286 VGND VPWR _0408_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[3\]
+ _0065_ sg13g2_dfrbpq_1
XFILLER_45_970 VPWR VGND sg13g2_decap_8
X_3931_ videogen.test_lut_thingy.pixel_feeder_inst.row\[22\]\[0\] net559 _1599_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_44_480 VPWR VGND sg13g2_decap_8
X_5100__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_20_815 VPWR VGND sg13g2_decap_4
X_3862_ net616 VPWR _1531_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[42\]\[3\]
+ net557 sg13g2_o21ai_1
XFILLER_32_653 VPWR VGND sg13g2_fill_1
X_2813_ net785 videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[0\] _0754_ _0493_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_859 VPWR VGND sg13g2_fill_2
X_3793_ _1461_ VPWR _1462_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[1\]
+ net586 sg13g2_o21ai_1
XFILLER_9_882 VPWR VGND sg13g2_decap_8
X_2744_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[1\] net777 _0738_ _0555_
+ VPWR VGND sg13g2_mux2_1
X_2675_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[1\] net773 _0717_ _0603_
+ VPWR VGND sg13g2_mux2_1
X_4414_ tmds_blue.dc_balancing_reg\[4\] _2056_ _2057_ VPWR VGND sg13g2_nor2_2
X_4345_ net606 _0862_ _1994_ VPWR VGND sg13g2_and2_1
XFILLER_28_1013 VPWR VGND sg13g2_decap_8
X_4276_ _1935_ _1934_ _1931_ _1938_ VPWR VGND sg13g2_a21o_1
X_3227_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[0\] _0940_ _0941_ VPWR VGND
+ sg13g2_and2_1
XFILLER_28_915 VPWR VGND sg13g2_decap_8
X_3158_ net548 _0886_ _0887_ VPWR VGND sg13g2_nor2_1
XFILLER_36_49 VPWR VGND sg13g2_decap_8
X_3089_ blue_tmds_par\[8\] net694 serialize.n429\[8\] VPWR VGND sg13g2_and2_1
XFILLER_14_119 VPWR VGND sg13g2_decap_4
XFILLER_35_480 VPWR VGND sg13g2_decap_8
XFILLER_11_815 VPWR VGND sg13g2_fill_1
XFILLER_11_848 VPWR VGND sg13g2_decap_4
XFILLER_10_347 VPWR VGND sg13g2_fill_2
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_46_767 VPWR VGND sg13g2_decap_4
XFILLER_18_458 VPWR VGND sg13g2_fill_2
XFILLER_27_970 VPWR VGND sg13g2_decap_8
XFILLER_34_929 VPWR VGND sg13g2_decap_8
XFILLER_26_491 VPWR VGND sg13g2_decap_4
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_10_881 VPWR VGND sg13g2_decap_8
XFILLER_6_852 VPWR VGND sg13g2_fill_1
X_4837__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_5_351 VPWR VGND sg13g2_fill_2
X_4130_ VGND VPWR _1794_ _1793_ _1791_ sg13g2_or2_1
XFILLER_3_42 VPWR VGND sg13g2_fill_1
X_4061_ _1724_ _1717_ _1713_ _1726_ VPWR VGND sg13g2_a21o_1
XFILLER_49_583 VPWR VGND sg13g2_decap_8
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
X_3012_ net746 videogen.test_lut_thingy.pixel_feeder_inst.state\[0\] _0808_ VPWR VGND
+ sg13g2_nor2_2
XFILLER_25_907 VPWR VGND sg13g2_decap_8
X_4963_ net319 VGND VPWR _0391_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[2\]
+ _0048_ sg13g2_dfrbpq_1
X_3914_ _1583_ net583 videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_33_973 VPWR VGND sg13g2_decap_8
X_4894_ net62 VGND VPWR _0322_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\]
+ net631 sg13g2_dfrbpq_2
XFILLER_20_634 VPWR VGND sg13g2_decap_4
X_3845_ videogen.test_lut_thingy.pixel_feeder_inst.row\[61\]\[3\] net563 _1514_ VPWR
+ VGND sg13g2_nor2_1
X_3776_ net612 _1433_ _1444_ _1445_ VPWR VGND sg13g2_nor3_1
X_2727_ net762 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\] _0734_ _0568_
+ VPWR VGND sg13g2_mux2_1
X_2658_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\] net773 _0708_ _0629_
+ VPWR VGND sg13g2_mux2_1
X_5031__182 VPWR VGND net182 sg13g2_tiehi
X_2589_ net614 _0645_ VPWR VGND sg13g2_inv_4
X_4328_ VGND VPWR _0914_ _1982_ _1984_ _1983_ sg13g2_a21oi_1
XFILLER_47_37 VPWR VGND sg13g2_decap_8
XFILLER_41_1021 VPWR VGND sg13g2_decap_8
X_4259_ _1921_ _1919_ _1920_ VPWR VGND sg13g2_nand2_1
XFILLER_27_200 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_15_406 VPWR VGND sg13g2_decap_4
XFILLER_24_962 VPWR VGND sg13g2_decap_8
XFILLER_11_612 VPWR VGND sg13g2_decap_8
XFILLER_23_461 VPWR VGND sg13g2_fill_2
XFILLER_11_656 VPWR VGND sg13g2_decap_8
XFILLER_10_155 VPWR VGND sg13g2_decap_4
XFILLER_11_678 VPWR VGND sg13g2_decap_8
XFILLER_3_822 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_2_343 VPWR VGND sg13g2_decap_4
XFILLER_3_899 VPWR VGND sg13g2_decap_8
Xfanout691 net692 net691 VPWR VGND sg13g2_buf_8
XFILLER_19_9 VPWR VGND sg13g2_decap_8
Xfanout680 net681 net680 VPWR VGND sg13g2_buf_8
XFILLER_34_726 VPWR VGND sg13g2_decap_8
XFILLER_15_940 VPWR VGND sg13g2_decap_8
XFILLER_30_910 VPWR VGND sg13g2_decap_8
X_5091__349 VPWR VGND net349 sg13g2_tiehi
X_3630_ _1296_ _1243_ _0662_ _1299_ VPWR VGND sg13g2_a21o_1
XFILLER_30_987 VPWR VGND sg13g2_decap_8
X_3561_ _1215_ _1211_ _1228_ _1230_ VPWR VGND sg13g2_a21o_1
X_3492_ _1103_ _1104_ _1101_ _1161_ VPWR VGND sg13g2_nand3_1
X_5231_ net800 VGND VPWR serialize.n429\[5\] serialize.n417\[3\] clknet_3_2__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5162_ net231 VGND VPWR _0586_ videogen.test_lut_thingy.pixel_feeder_inst.row\[1\]\[0\]
+ _0234_ sg13g2_dfrbpq_1
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
X_5093_ net318 VGND VPWR _0517_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[3\]
+ _0165_ sg13g2_dfrbpq_1
X_4113_ _1777_ _1703_ _1778_ VPWR VGND sg13g2_xor2_1
X_4044_ _1093_ _1706_ _1709_ VPWR VGND sg13g2_nor2_1
XFILLER_37_586 VPWR VGND sg13g2_decap_8
XFILLER_24_203 VPWR VGND sg13g2_decap_4
XFILLER_24_236 VPWR VGND sg13g2_fill_2
XFILLER_25_759 VPWR VGND sg13g2_decap_8
XFILLER_24_269 VPWR VGND sg13g2_fill_1
X_4946_ net338 VGND VPWR _0374_ tmds_blue.n126 net636 sg13g2_dfrbpq_1
X_4877_ net91 VGND VPWR _0305_ videogen.fancy_shader.video_x\[6\] net634 sg13g2_dfrbpq_2
XFILLER_21_943 VPWR VGND sg13g2_decap_8
X_3828_ net615 VPWR _1497_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[56\]\[3\]
+ net586 sg13g2_o21ai_1
XFILLER_20_453 VPWR VGND sg13g2_fill_1
X_3759_ net618 VPWR _1428_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[1\]
+ net550 sg13g2_o21ai_1
XFILLER_3_118 VPWR VGND sg13g2_decap_8
XFILLER_0_803 VPWR VGND sg13g2_decap_8
X_5183__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_28_553 VPWR VGND sg13g2_fill_2
XFILLER_15_236 VPWR VGND sg13g2_fill_1
XFILLER_11_442 VPWR VGND sg13g2_fill_2
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_8_947 VPWR VGND sg13g2_decap_8
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_674 VPWR VGND sg13g2_fill_1
XFILLER_2_195 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_fill_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_46_394 VPWR VGND sg13g2_fill_2
XFILLER_46_383 VPWR VGND sg13g2_decap_8
XFILLER_34_534 VPWR VGND sg13g2_decap_4
X_4800_ net690 net741 _0230_ VPWR VGND sg13g2_nor2_1
X_5195__148 VPWR VGND net148 sg13g2_tiehi
X_2992_ _0707_ _0714_ _0801_ VPWR VGND sg13g2_nor2_2
X_4731_ net650 net702 _0161_ VPWR VGND sg13g2_nor2_1
X_4662_ net684 net736 _0092_ VPWR VGND sg13g2_nor2_1
X_3613_ _1282_ _1066_ _1279_ VPWR VGND sg13g2_xnor2_1
X_4593_ net649 net701 _0023_ VPWR VGND sg13g2_nor2_1
X_3544_ _1208_ _1212_ _1213_ VPWR VGND sg13g2_and2_1
X_3475_ _1094_ _1095_ _1099_ _1144_ VPWR VGND sg13g2_or3_1
X_5214_ net801 VGND VPWR serialize.n428\[6\] serialize.n414\[4\] clknet_3_4__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_5145_ net37 VGND VPWR _0569_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\]
+ _0217_ sg13g2_dfrbpq_1
X_5076_ net391 VGND VPWR _0500_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[3\]
+ _0157_ sg13g2_dfrbpq_1
X_4027_ _1695_ _1495_ _1693_ VPWR VGND sg13g2_nand2_1
XFILLER_25_534 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_fill_1
XFILLER_25_545 VPWR VGND sg13g2_decap_8
XFILLER_25_589 VPWR VGND sg13g2_decap_8
X_5000__243 VPWR VGND net243 sg13g2_tiehi
X_4929_ net364 VGND VPWR _0357_ videogen.fancy_shader.video_y\[1\] net633 sg13g2_dfrbpq_2
X_4857__125 VPWR VGND net125 sg13g2_tiehi
X_5074__399 VPWR VGND net399 sg13g2_tiehi
XFILLER_4_438 VPWR VGND sg13g2_decap_8
Xheichips25_bagel_21 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_0_655 VPWR VGND sg13g2_decap_4
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_47_125 VPWR VGND sg13g2_fill_2
XFILLER_47_114 VPWR VGND sg13g2_decap_8
X_5069__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_28_350 VPWR VGND sg13g2_decap_4
XFILLER_29_851 VPWR VGND sg13g2_decap_8
XFILLER_29_895 VPWR VGND sg13g2_fill_2
XFILLER_43_353 VPWR VGND sg13g2_fill_1
XFILLER_43_342 VPWR VGND sg13g2_decap_8
XFILLER_16_589 VPWR VGND sg13g2_decap_4
X_4840__151 VPWR VGND net151 sg13g2_tiehi
XFILLER_8_700 VPWR VGND sg13g2_decap_8
XFILLER_12_762 VPWR VGND sg13g2_decap_8
XFILLER_11_272 VPWR VGND sg13g2_fill_1
XFILLER_8_788 VPWR VGND sg13g2_decap_8
X_3260_ VGND VPWR _0964_ _0963_ net611 sg13g2_or2_1
XFILLER_38_103 VPWR VGND sg13g2_fill_1
X_3191_ _0852_ VPWR _0918_ VGND _0882_ _0917_ sg13g2_o21ai_1
XFILLER_39_659 VPWR VGND sg13g2_decap_8
XFILLER_35_832 VPWR VGND sg13g2_fill_2
XFILLER_34_331 VPWR VGND sg13g2_decap_8
XFILLER_34_364 VPWR VGND sg13g2_decap_8
XFILLER_14_19 VPWR VGND sg13g2_fill_1
XFILLER_34_397 VPWR VGND sg13g2_fill_1
X_4714_ net674 net726 _0144_ VPWR VGND sg13g2_nor2_1
X_2975_ _0796_ _0716_ _0781_ VPWR VGND sg13g2_nand2_2
X_4645_ net669 net722 _0075_ VPWR VGND sg13g2_nor2_1
X_4576_ net674 net726 _0008_ VPWR VGND sg13g2_nor2_1
X_3527_ _1196_ _1193_ _1194_ VPWR VGND sg13g2_nand2_1
XFILLER_39_27 VPWR VGND sg13g2_decap_8
X_3458_ _1124_ _1122_ _1125_ _1127_ VPWR VGND sg13g2_a21o_2
X_3389_ VGND VPWR _1057_ _1058_ _0370_ net745 sg13g2_a21oi_1
XFILLER_29_125 VPWR VGND sg13g2_fill_1
X_5128_ net177 VGND VPWR _0552_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[2\]
+ _0200_ sg13g2_dfrbpq_1
XFILLER_29_158 VPWR VGND sg13g2_decap_4
X_5059_ net72 VGND VPWR _0487_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[2\]
+ _0144_ sg13g2_dfrbpq_1
XFILLER_26_832 VPWR VGND sg13g2_decap_8
XFILLER_25_342 VPWR VGND sg13g2_decap_4
XFILLER_13_526 VPWR VGND sg13g2_decap_4
XFILLER_40_378 VPWR VGND sg13g2_decap_4
XFILLER_40_367 VPWR VGND sg13g2_decap_8
XFILLER_21_592 VPWR VGND sg13g2_decap_8
XFILLER_45_1019 VPWR VGND sg13g2_decap_4
XFILLER_1_942 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_48_401 VPWR VGND sg13g2_decap_4
XFILLER_0_474 VPWR VGND sg13g2_decap_8
XFILLER_29_71 VPWR VGND sg13g2_fill_1
XFILLER_44_651 VPWR VGND sg13g2_fill_1
XFILLER_45_92 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_fill_2
XFILLER_17_898 VPWR VGND sg13g2_decap_8
XFILLER_43_194 VPWR VGND sg13g2_decap_8
XFILLER_32_857 VPWR VGND sg13g2_fill_2
X_2760_ videogen.test_lut_thingy.pixel_feeder_inst.row\[30\]\[0\] net788 _0741_ _0542_
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_541 VPWR VGND sg13g2_fill_2
X_2691_ _0712_ _0719_ _0724_ VPWR VGND sg13g2_nor2_2
X_4430_ VGND VPWR net603 _2057_ _2070_ _2061_ sg13g2_a21oi_1
X_4361_ VPWR _2007_ _2006_ VGND sg13g2_inv_1
X_3312_ videogen.fancy_shader.video_x\[2\] videogen.fancy_shader.n646\[2\] _1002_
+ VPWR VGND sg13g2_xor2_1
X_4292_ VGND VPWR _1950_ _1953_ _1954_ _1948_ sg13g2_a21oi_1
X_3243_ _0943_ _0951_ _0952_ _0322_ VPWR VGND sg13g2_nor3_1
X_3174_ _0901_ _0902_ _0903_ VPWR VGND sg13g2_nor2_1
XFILLER_35_640 VPWR VGND sg13g2_fill_2
XFILLER_23_813 VPWR VGND sg13g2_decap_8
X_2958_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[1\] net782 _0792_ _0343_
+ VPWR VGND sg13g2_mux2_1
X_2889_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[1\] _0775_ _0438_
+ VPWR VGND sg13g2_mux2_1
X_4628_ net652 net704 _0058_ VPWR VGND sg13g2_nor2_1
X_4559_ VGND VPWR _2134_ _2156_ _2188_ _2187_ sg13g2_a21oi_1
XFILLER_46_916 VPWR VGND sg13g2_decap_8
XFILLER_39_990 VPWR VGND sg13g2_decap_8
X_5041__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_9_338 VPWR VGND sg13g2_fill_1
Xoutput4 net4 tmds_clk VPWR VGND sg13g2_buf_1
XFILLER_5_599 VPWR VGND sg13g2_fill_2
XFILLER_0_260 VPWR VGND sg13g2_decap_8
XFILLER_49_798 VPWR VGND sg13g2_decap_8
XFILLER_36_448 VPWR VGND sg13g2_decap_4
X_3930_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[0\] net591 _1598_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_44_470 VPWR VGND sg13g2_decap_4
X_5094__314 VPWR VGND net314 sg13g2_tiehi
XFILLER_32_632 VPWR VGND sg13g2_decap_8
X_3861_ videogen.test_lut_thingy.pixel_feeder_inst.row\[43\]\[3\] net579 _1530_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_31_131 VPWR VGND sg13g2_decap_8
X_3792_ VGND VPWR _1461_ net563 videogen.test_lut_thingy.pixel_feeder_inst.row\[57\]\[1\]
+ sg13g2_or2_1
X_2812_ net774 videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[1\] _0754_ _0494_
+ VPWR VGND sg13g2_mux2_1
XFILLER_20_827 VPWR VGND sg13g2_decap_8
X_2743_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[2\] net769 _0738_ _0556_
+ VPWR VGND sg13g2_mux2_1
X_2674_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[2\] net762 _0717_ _0604_
+ VPWR VGND sg13g2_mux2_1
X_4413_ tmds_blue.dc_balancing_reg\[0\] tmds_blue.dc_balancing_reg\[1\] tmds_blue.dc_balancing_reg\[3\]
+ tmds_blue.dc_balancing_reg\[2\] _2056_ VPWR VGND sg13g2_or4_1
X_4344_ VGND VPWR tmds_green.n100 net605 _0507_ net749 sg13g2_a21oi_1
X_4275_ VGND VPWR _1934_ _1935_ _1937_ _1931_ sg13g2_a21oi_1
XFILLER_39_253 VPWR VGND sg13g2_decap_8
X_3226_ _0938_ _0939_ _0940_ VPWR VGND sg13g2_nor2_2
X_3157_ tmds_red.n102 _0885_ _0886_ VPWR VGND sg13g2_nor2_1
X_3088_ net425 blue_tmds_par\[7\] net694 serialize.n429\[7\] VPWR VGND sg13g2_mux2_1
XFILLER_42_407 VPWR VGND sg13g2_decap_4
XFILLER_23_665 VPWR VGND sg13g2_fill_1
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_fill_1
XFILLER_10_359 VPWR VGND sg13g2_decap_8
X_4975__296 VPWR VGND net296 sg13g2_tiehi
XFILLER_19_916 VPWR VGND sg13g2_decap_8
XFILLER_34_908 VPWR VGND sg13g2_decap_8
XFILLER_33_407 VPWR VGND sg13g2_fill_2
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_26_72 VPWR VGND sg13g2_fill_1
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_13_142 VPWR VGND sg13g2_decap_8
XFILLER_9_113 VPWR VGND sg13g2_fill_2
XFILLER_13_153 VPWR VGND sg13g2_fill_2
XFILLER_14_676 VPWR VGND sg13g2_fill_1
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_3_65 VPWR VGND sg13g2_decap_8
X_4060_ _1718_ _1719_ _1721_ _1722_ _1725_ VPWR VGND sg13g2_or4_1
XFILLER_3_98 VPWR VGND sg13g2_fill_2
XFILLER_49_562 VPWR VGND sg13g2_decap_8
X_3011_ net795 _0807_ _0371_ VPWR VGND sg13g2_and2_1
XFILLER_37_768 VPWR VGND sg13g2_decap_8
XFILLER_37_757 VPWR VGND sg13g2_fill_1
XFILLER_18_982 VPWR VGND sg13g2_decap_8
X_4962_ net321 VGND VPWR _0390_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[1\]
+ _0047_ sg13g2_dfrbpq_1
X_4893_ net64 VGND VPWR _0321_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[3\]
+ net631 sg13g2_dfrbpq_2
X_3913_ videogen.test_lut_thingy.pixel_feeder_inst.row\[26\]\[3\] net552 _1582_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_32_451 VPWR VGND sg13g2_fill_2
XFILLER_33_952 VPWR VGND sg13g2_decap_8
X_3844_ net615 VPWR _1513_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[3\]
+ net553 sg13g2_o21ai_1
XFILLER_22_19 VPWR VGND sg13g2_fill_1
X_3775_ net614 _1438_ _1443_ _1444_ VPWR VGND sg13g2_nor3_1
X_2726_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[3\] _0734_ _0569_
+ VPWR VGND sg13g2_mux2_1
X_2657_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[2\] net763 _0708_ _0630_
+ VPWR VGND sg13g2_mux2_1
X_2588_ VPWR _0644_ net611 VGND sg13g2_inv_1
X_4327_ net606 VPWR _1983_ VGND _0914_ _1982_ sg13g2_o21ai_1
XFILLER_41_1000 VPWR VGND sg13g2_decap_8
X_4258_ _1903_ _1910_ _1918_ _1920_ VPWR VGND sg13g2_or3_1
X_3209_ _0815_ _0923_ _0928_ _0304_ VPWR VGND sg13g2_nor3_1
X_4189_ _1851_ _1827_ _1850_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_705 VPWR VGND sg13g2_fill_1
XFILLER_42_215 VPWR VGND sg13g2_decap_8
XFILLER_42_248 VPWR VGND sg13g2_decap_8
XFILLER_23_440 VPWR VGND sg13g2_decap_4
XFILLER_24_941 VPWR VGND sg13g2_decap_8
XFILLER_12_41 VPWR VGND sg13g2_fill_1
XFILLER_3_801 VPWR VGND sg13g2_decap_8
XFILLER_5_2 VPWR VGND sg13g2_fill_1
XFILLER_3_878 VPWR VGND sg13g2_decap_8
XFILLER_2_366 VPWR VGND sg13g2_fill_2
X_4867__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_2_399 VPWR VGND sg13g2_decap_8
Xfanout692 net693 net692 VPWR VGND sg13g2_buf_2
Xfanout670 net671 net670 VPWR VGND sg13g2_buf_8
Xfanout681 net682 net681 VPWR VGND sg13g2_buf_2
XFILLER_46_521 VPWR VGND sg13g2_fill_1
XFILLER_37_82 VPWR VGND sg13g2_decap_8
XFILLER_18_245 VPWR VGND sg13g2_decap_8
XFILLER_34_705 VPWR VGND sg13g2_decap_8
XFILLER_14_462 VPWR VGND sg13g2_fill_2
XFILLER_15_996 VPWR VGND sg13g2_decap_8
XFILLER_18_1024 VPWR VGND sg13g2_decap_4
XFILLER_14_495 VPWR VGND sg13g2_decap_8
XFILLER_30_966 VPWR VGND sg13g2_decap_8
X_3560_ VGND VPWR _1211_ _1215_ _1229_ _1228_ sg13g2_a21oi_1
X_5230_ net800 VGND VPWR net444 serialize.n417\[2\] clknet_3_1__leaf_clk_regs sg13g2_dfrbpq_1
X_3491_ _1160_ _1127_ _1159_ VPWR VGND sg13g2_nand2_1
X_5161_ net238 VGND VPWR _0585_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[3\]
+ _0233_ sg13g2_dfrbpq_1
X_5092_ net322 VGND VPWR _0516_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[2\]
+ _0164_ sg13g2_dfrbpq_1
X_4112_ VGND VPWR _1767_ _1777_ _1776_ _1772_ sg13g2_a21oi_2
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4043_ _1073_ _1706_ _1708_ VPWR VGND sg13g2_nor2_1
XFILLER_25_749 VPWR VGND sg13g2_decap_4
X_4945_ net339 VGND VPWR _0373_ tmds_blue.n100 net636 sg13g2_dfrbpq_1
XFILLER_21_922 VPWR VGND sg13g2_decap_8
X_4876_ net92 VGND VPWR _0304_ videogen.fancy_shader.video_x\[5\] net634 sg13g2_dfrbpq_2
XFILLER_32_281 VPWR VGND sg13g2_fill_2
XFILLER_20_465 VPWR VGND sg13g2_decap_8
XFILLER_20_476 VPWR VGND sg13g2_fill_1
XFILLER_21_999 VPWR VGND sg13g2_decap_8
X_3827_ _1399_ _1495_ _1496_ VPWR VGND sg13g2_nor2_1
X_3758_ net618 _1423_ _1424_ _1426_ _1427_ VPWR VGND sg13g2_nor4_1
X_2709_ videogen.test_lut_thingy.pixel_feeder_inst.row\[21\]\[3\] net760 _0729_ _0581_
+ VPWR VGND sg13g2_mux2_1
X_3689_ videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\] net558 _1358_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_0_859 VPWR VGND sg13g2_decap_8
XFILLER_28_510 VPWR VGND sg13g2_decap_8
XFILLER_43_513 VPWR VGND sg13g2_fill_1
XFILLER_28_587 VPWR VGND sg13g2_decap_4
XFILLER_31_708 VPWR VGND sg13g2_fill_1
XFILLER_12_933 VPWR VGND sg13g2_decap_8
XFILLER_8_926 VPWR VGND sg13g2_decap_8
XFILLER_11_454 VPWR VGND sg13g2_fill_2
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_808 VPWR VGND sg13g2_fill_1
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_46_351 VPWR VGND sg13g2_decap_4
XFILLER_19_565 VPWR VGND sg13g2_decap_4
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_46_373 VPWR VGND sg13g2_decap_4
XFILLER_0_55 VPWR VGND sg13g2_fill_1
XFILLER_19_587 VPWR VGND sg13g2_decap_8
XFILLER_34_546 VPWR VGND sg13g2_fill_2
X_2991_ net791 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\] _0800_ _0287_
+ VPWR VGND sg13g2_mux2_1
X_4730_ net650 net702 _0160_ VPWR VGND sg13g2_nor2_1
X_4661_ net684 net736 _0091_ VPWR VGND sg13g2_nor2_1
XFILLER_30_774 VPWR VGND sg13g2_decap_8
X_3612_ _1281_ _1267_ _1280_ VPWR VGND sg13g2_xnor2_1
X_4592_ net649 net701 _0022_ VPWR VGND sg13g2_nor2_1
X_3543_ _1201_ _1205_ _1195_ _1212_ VPWR VGND sg13g2_nand3_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_3474_ _1099_ VPWR _1143_ VGND _1094_ _1095_ sg13g2_o21ai_1
X_5213_ net803 VGND VPWR serialize.n428\[5\] serialize.n414\[3\] clknet_3_6__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
X_5144_ net45 VGND VPWR _0568_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[2\]
+ _0216_ sg13g2_dfrbpq_1
XFILLER_29_318 VPWR VGND sg13g2_decap_8
X_5075_ net395 VGND VPWR _0499_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[2\]
+ _0156_ sg13g2_dfrbpq_1
XFILLER_38_874 VPWR VGND sg13g2_decap_8
XFILLER_37_340 VPWR VGND sg13g2_decap_8
X_4026_ VPWR _1694_ _1693_ VGND sg13g2_inv_1
XFILLER_13_708 VPWR VGND sg13g2_fill_1
XFILLER_40_505 VPWR VGND sg13g2_fill_1
XFILLER_12_229 VPWR VGND sg13g2_decap_8
X_4928_ net366 VGND VPWR _0356_ videogen.fancy_shader.video_y\[0\] net633 sg13g2_dfrbpq_1
XFILLER_21_774 VPWR VGND sg13g2_fill_2
X_4859_ net121 VGND VPWR _0287_ videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[0\]
+ _0018_ sg13g2_dfrbpq_1
Xheichips25_bagel_22 VPWR VGND uio_oe[3] sg13g2_tielo
XFILLER_48_638 VPWR VGND sg13g2_fill_1
XFILLER_47_148 VPWR VGND sg13g2_decap_4
XFILLER_18_51 VPWR VGND sg13g2_fill_2
XFILLER_44_844 VPWR VGND sg13g2_decap_8
XFILLER_16_546 VPWR VGND sg13g2_decap_8
XFILLER_24_590 VPWR VGND sg13g2_decap_8
XFILLER_34_72 VPWR VGND sg13g2_decap_8
XFILLER_8_734 VPWR VGND sg13g2_fill_1
XFILLER_8_778 VPWR VGND sg13g2_fill_2
XFILLER_4_995 VPWR VGND sg13g2_decap_8
XFILLER_3_461 VPWR VGND sg13g2_fill_2
XFILLER_39_605 VPWR VGND sg13g2_decap_8
X_3190_ net571 _0917_ _0275_ VPWR VGND sg13g2_nor2_1
XFILLER_38_115 VPWR VGND sg13g2_decap_4
XFILLER_15_4 VPWR VGND sg13g2_decap_4
XFILLER_22_1009 VPWR VGND sg13g2_decap_8
XFILLER_38_148 VPWR VGND sg13g2_decap_4
XFILLER_19_384 VPWR VGND sg13g2_fill_2
XFILLER_22_505 VPWR VGND sg13g2_decap_8
XFILLER_22_527 VPWR VGND sg13g2_decap_4
X_2974_ net786 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[0\] _0795_ _0309_
+ VPWR VGND sg13g2_mux2_1
X_4713_ net677 net726 _0143_ VPWR VGND sg13g2_nor2_1
X_4644_ net669 net722 _0074_ VPWR VGND sg13g2_nor2_1
X_4575_ net674 net726 _0007_ VPWR VGND sg13g2_nor2_1
X_3526_ _1193_ _1194_ _1195_ VPWR VGND sg13g2_and2_1
X_3457_ VGND VPWR _1122_ _1124_ _1126_ _1125_ sg13g2_a21oi_1
X_3388_ VGND VPWR _0678_ _0813_ _1058_ _0805_ sg13g2_a21oi_1
XFILLER_29_115 VPWR VGND sg13g2_fill_1
X_5127_ net181 VGND VPWR _0551_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[1\]
+ _0199_ sg13g2_dfrbpq_1
X_5058_ net76 VGND VPWR _0486_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[1\]
+ _0143_ sg13g2_dfrbpq_1
X_5028__188 VPWR VGND net188 sg13g2_tiehi
X_4009_ _1673_ _1674_ _1675_ _1676_ _1677_ VPWR VGND sg13g2_nor4_1
XFILLER_26_811 VPWR VGND sg13g2_decap_8
XFILLER_41_814 VPWR VGND sg13g2_decap_8
XFILLER_13_505 VPWR VGND sg13g2_decap_8
XFILLER_25_376 VPWR VGND sg13g2_fill_2
XFILLER_26_888 VPWR VGND sg13g2_decap_8
XFILLER_40_313 VPWR VGND sg13g2_decap_8
XFILLER_1_921 VPWR VGND sg13g2_decap_8
X_4888__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_49_903 VPWR VGND sg13g2_decap_8
XFILLER_0_453 VPWR VGND sg13g2_decap_8
X_4985__276 VPWR VGND net276 sg13g2_tiehi
XFILLER_1_998 VPWR VGND sg13g2_decap_8
XFILLER_21_1020 VPWR VGND sg13g2_decap_8
XFILLER_29_83 VPWR VGND sg13g2_fill_1
XFILLER_45_60 VPWR VGND sg13g2_fill_2
XFILLER_16_387 VPWR VGND sg13g2_fill_2
XFILLER_8_520 VPWR VGND sg13g2_decap_8
X_2690_ net792 videogen.test_lut_thingy.pixel_feeder_inst.row\[17\]\[0\] _0723_ _0594_
+ VPWR VGND sg13g2_mux2_1
X_4360_ net547 _2005_ _2006_ VPWR VGND sg13g2_nor2_1
X_3311_ videogen.fancy_shader.n646\[2\] videogen.fancy_shader.video_x\[2\] _1001_
+ VPWR VGND sg13g2_and2_1
X_4291_ _1953_ _1951_ _1952_ VPWR VGND sg13g2_xnor2_1
X_3242_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0950_ _0952_ VPWR VGND
+ sg13g2_and2_1
X_3173_ _0899_ _0900_ _0902_ VPWR VGND sg13g2_nor2b_2
XFILLER_48_991 VPWR VGND sg13g2_decap_8
XFILLER_19_170 VPWR VGND sg13g2_fill_1
X_5056__84 VPWR VGND net84 sg13g2_tiehi
XFILLER_35_674 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_4
XFILLER_22_357 VPWR VGND sg13g2_decap_4
XFILLER_31_880 VPWR VGND sg13g2_fill_1
X_2957_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[2\] net770 _0792_ _0344_
+ VPWR VGND sg13g2_mux2_1
X_2888_ net771 videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[2\] _0775_ _0439_
+ VPWR VGND sg13g2_mux2_1
X_4627_ net663 net713 _0057_ VPWR VGND sg13g2_nor2_1
X_4558_ _2170_ _2186_ _2187_ VPWR VGND sg13g2_nor2b_1
X_4489_ _2109_ _2121_ _2122_ VPWR VGND sg13g2_nor2_1
X_3509_ _1178_ net544 _1176_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_1020 VPWR VGND sg13g2_decap_8
X_5141__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_41_600 VPWR VGND sg13g2_decap_8
XFILLER_13_313 VPWR VGND sg13g2_decap_4
XFILLER_14_825 VPWR VGND sg13g2_decap_8
XFILLER_13_357 VPWR VGND sg13g2_fill_1
XFILLER_40_176 VPWR VGND sg13g2_decap_8
XFILLER_13_379 VPWR VGND sg13g2_fill_2
XFILLER_31_84 VPWR VGND sg13g2_decap_8
XFILLER_5_578 VPWR VGND sg13g2_decap_8
Xoutput5 net5 tmds_g VPWR VGND sg13g2_buf_1
XFILLER_1_795 VPWR VGND sg13g2_decap_8
XFILLER_49_766 VPWR VGND sg13g2_decap_4
XFILLER_37_906 VPWR VGND sg13g2_fill_1
X_4891__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_16_162 VPWR VGND sg13g2_fill_2
XFILLER_32_611 VPWR VGND sg13g2_decap_8
X_3860_ videogen.test_lut_thingy.pixel_feeder_inst.row\[40\]\[3\] net589 _1529_ VPWR
+ VGND sg13g2_nor2_1
X_3791_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[1\] net575 _1460_ VPWR
+ VGND sg13g2_nor2_1
X_2811_ net763 videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[2\] _0754_ _0495_
+ VPWR VGND sg13g2_mux2_1
XFILLER_31_165 VPWR VGND sg13g2_fill_2
XFILLER_13_891 VPWR VGND sg13g2_decap_8
X_2742_ videogen.test_lut_thingy.pixel_feeder_inst.row\[27\]\[3\] net752 _0738_ _0557_
+ VPWR VGND sg13g2_mux2_1
X_2673_ videogen.test_lut_thingy.pixel_feeder_inst.row\[7\]\[3\] net753 _0717_ _0605_
+ VPWR VGND sg13g2_mux2_1
X_4412_ VGND VPWR _2054_ _2055_ _0513_ net572 sg13g2_a21oi_1
X_4343_ net748 _1993_ _0506_ VPWR VGND sg13g2_nor2_1
X_4274_ _1936_ _1934_ _1935_ VPWR VGND sg13g2_nand2_1
X_3225_ _0684_ VPWR _0939_ VGND videogen.test_lut_thingy.pixel_feeder_inst.state\[2\]
+ _0824_ sg13g2_o21ai_1
XFILLER_39_232 VPWR VGND sg13g2_fill_1
X_3156_ _0885_ _0869_ _0883_ VPWR VGND sg13g2_xnor2_1
X_3087_ net435 blue_tmds_par\[6\] net694 serialize.n429\[6\] VPWR VGND sg13g2_mux2_1
XFILLER_39_298 VPWR VGND sg13g2_fill_2
XFILLER_36_983 VPWR VGND sg13g2_decap_8
XFILLER_23_633 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_fill_1
X_3989_ videogen.test_lut_thingy.pixel_feeder_inst.row\[59\]\[0\] net576 _1657_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_10_349 VPWR VGND sg13g2_fill_1
XFILLER_45_235 VPWR VGND sg13g2_decap_8
XFILLER_14_622 VPWR VGND sg13g2_decap_8
XFILLER_9_125 VPWR VGND sg13g2_decap_8
XFILLER_9_136 VPWR VGND sg13g2_fill_2
XFILLER_6_843 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_33 VPWR VGND sg13g2_fill_1
XFILLER_49_541 VPWR VGND sg13g2_decap_8
X_3010_ videogen.fancy_shader.video_y\[9\] _0674_ _0804_ _0807_ VGND VPWR _0806_ sg13g2_nor4_2
XFILLER_36_224 VPWR VGND sg13g2_fill_2
XFILLER_18_961 VPWR VGND sg13g2_decap_8
X_4961_ net323 VGND VPWR _0389_ videogen.test_lut_thingy.pixel_feeder_inst.row\[62\]\[0\]
+ _0046_ sg13g2_dfrbpq_1
XFILLER_33_931 VPWR VGND sg13g2_decap_8
X_4892_ net66 VGND VPWR _0320_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[2\]
+ net631 sg13g2_dfrbpq_2
X_3912_ _1577_ _1578_ _1579_ _1580_ _1581_ VPWR VGND sg13g2_nor4_1
X_3843_ _1508_ _1509_ _1510_ _1511_ _1512_ VPWR VGND sg13g2_nor4_1
XFILLER_9_670 VPWR VGND sg13g2_fill_2
X_3774_ net621 _1439_ _1440_ _1442_ _1443_ VPWR VGND sg13g2_nor4_1
X_2725_ _0734_ _0720_ _0732_ VPWR VGND sg13g2_nand2_2
X_2656_ videogen.test_lut_thingy.pixel_feeder_inst.row\[14\]\[3\] net753 _0708_ _0631_
+ VPWR VGND sg13g2_mux2_1
X_2587_ VPWR _0643_ videogen.fancy_shader.n646\[0\] VGND sg13g2_inv_1
X_4326_ _0882_ tmds_red.n114 _1982_ VPWR VGND sg13g2_xor2_1
XFILLER_47_28 VPWR VGND sg13g2_decap_4
X_4257_ _1918_ VPWR _1919_ VGND _1903_ _1910_ sg13g2_o21ai_1
X_3208_ videogen.fancy_shader.video_x\[5\] _0814_ _0928_ VPWR VGND sg13g2_nor2_1
X_4188_ _1837_ VPWR _1850_ VGND _1847_ _1849_ sg13g2_o21ai_1
X_3139_ tmds_red.n114 tmds_red.n132 _0868_ VPWR VGND sg13g2_nor2_1
XFILLER_28_736 VPWR VGND sg13g2_decap_4
XFILLER_24_920 VPWR VGND sg13g2_decap_8
XFILLER_24_997 VPWR VGND sg13g2_decap_8
XFILLER_10_113 VPWR VGND sg13g2_fill_1
X_5077__387 VPWR VGND net387 sg13g2_tiehi
XFILLER_10_168 VPWR VGND sg13g2_decap_4
XFILLER_6_128 VPWR VGND sg13g2_decap_8
X_5010__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xfanout660 net662 net660 VPWR VGND sg13g2_buf_8
Xfanout693 clockdiv.q2temp net693 VPWR VGND sg13g2_buf_8
Xfanout682 net693 net682 VPWR VGND sg13g2_buf_8
Xfanout671 net672 net671 VPWR VGND sg13g2_buf_8
X_5160__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_18_235 VPWR VGND sg13g2_decap_4
XFILLER_18_257 VPWR VGND sg13g2_decap_8
XFILLER_18_268 VPWR VGND sg13g2_fill_1
XFILLER_27_780 VPWR VGND sg13g2_fill_1
XFILLER_18_1003 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_decap_8
XFILLER_33_249 VPWR VGND sg13g2_fill_2
XFILLER_15_975 VPWR VGND sg13g2_decap_8
XFILLER_30_945 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk_regs clknet_0_clk_regs clknet_3_7__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_6_662 VPWR VGND sg13g2_fill_1
X_3490_ _1124_ _1125_ _1122_ _1159_ VPWR VGND sg13g2_nand3_1
XFILLER_6_684 VPWR VGND sg13g2_decap_4
XFILLER_5_150 VPWR VGND sg13g2_fill_2
X_5160_ net246 VGND VPWR _0584_ videogen.test_lut_thingy.pixel_feeder_inst.row\[20\]\[2\]
+ _0232_ sg13g2_dfrbpq_1
X_5091_ net349 VGND VPWR _0515_ videogen.test_lut_thingy.pixel_feeder_inst.row\[37\]\[1\]
+ _0163_ sg13g2_dfrbpq_1
X_4111_ _1776_ _1773_ _1775_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_360 VPWR VGND sg13g2_decap_8
X_4042_ _1707_ _1076_ _1706_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_371 VPWR VGND sg13g2_fill_1
XFILLER_37_577 VPWR VGND sg13g2_fill_1
XFILLER_18_780 VPWR VGND sg13g2_decap_4
X_4944_ net340 VGND VPWR _0372_ tmds_blue.n193 net636 sg13g2_dfrbpq_2
XFILLER_21_901 VPWR VGND sg13g2_decap_8
XFILLER_33_783 VPWR VGND sg13g2_decap_8
X_4875_ net93 VGND VPWR _0303_ videogen.fancy_shader.video_x\[4\] net633 sg13g2_dfrbpq_2
XFILLER_20_411 VPWR VGND sg13g2_decap_8
XFILLER_32_293 VPWR VGND sg13g2_fill_1
XFILLER_21_978 VPWR VGND sg13g2_decap_8
X_3826_ _1494_ VPWR _1495_ VGND _0660_ net2 sg13g2_o21ai_1
X_3757_ _1425_ VPWR _1426_ VGND videogen.test_lut_thingy.pixel_feeder_inst.row\[10\]\[1\]
+ net550 sg13g2_o21ai_1
X_2708_ _0719_ _0728_ _0729_ VPWR VGND sg13g2_nor2_2
X_3688_ videogen.test_lut_thingy.pixel_feeder_inst.row\[48\]\[2\] net590 _1357_ VPWR
+ VGND sg13g2_nor2_1
X_2639_ _0644_ _0689_ _0692_ VPWR VGND sg13g2_and2_1
XFILLER_0_838 VPWR VGND sg13g2_decap_8
X_4309_ VPWR VGND _1961_ _1970_ _1966_ _1857_ _1971_ _1965_ sg13g2_a221oi_1
XFILLER_28_566 VPWR VGND sg13g2_decap_8
XFILLER_43_569 VPWR VGND sg13g2_fill_2
XFILLER_15_227 VPWR VGND sg13g2_fill_2
XFILLER_12_912 VPWR VGND sg13g2_decap_8
XFILLER_24_772 VPWR VGND sg13g2_decap_4
XFILLER_8_905 VPWR VGND sg13g2_decap_8
XFILLER_23_282 VPWR VGND sg13g2_fill_2
XFILLER_12_989 VPWR VGND sg13g2_decap_8
X_5038__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_23_293 VPWR VGND sg13g2_decap_8
XFILLER_3_632 VPWR VGND sg13g2_decap_8
XFILLER_3_698 VPWR VGND sg13g2_decap_4
XFILLER_2_142 VPWR VGND sg13g2_decap_8
XFILLER_24_9 VPWR VGND sg13g2_decap_8
XFILLER_47_831 VPWR VGND sg13g2_fill_2
XFILLER_47_820 VPWR VGND sg13g2_decap_8
XFILLER_19_500 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_fill_1
XFILLER_19_522 VPWR VGND sg13g2_fill_2
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_46_341 VPWR VGND sg13g2_fill_1
XFILLER_46_330 VPWR VGND sg13g2_decap_8
XFILLER_0_67 VPWR VGND sg13g2_decap_8
X_2990_ net781 videogen.test_lut_thingy.pixel_feeder_inst.row\[49\]\[1\] _0800_ _0288_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_772 VPWR VGND sg13g2_decap_4
X_4660_ net684 net736 _0090_ VPWR VGND sg13g2_nor2_1
XFILLER_30_742 VPWR VGND sg13g2_fill_1
X_3611_ VGND VPWR _1276_ _1279_ _1280_ _1273_ sg13g2_a21oi_1
X_4591_ net684 net736 _0021_ VPWR VGND sg13g2_nor2_1
XFILLER_6_470 VPWR VGND sg13g2_fill_1
X_3542_ _1207_ VPWR _1211_ VGND _1209_ _1210_ sg13g2_o21ai_1
X_3473_ _1140_ _1141_ _1142_ VPWR VGND sg13g2_and2_1
X_5212_ net802 VGND VPWR serialize.n428\[4\] serialize.n414\[2\] clknet_3_5__leaf_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
X_5143_ net53 VGND VPWR _0567_ videogen.test_lut_thingy.pixel_feeder_inst.row\[24\]\[1\]
+ _0215_ sg13g2_dfrbpq_1
XFILLER_36_0 VPWR VGND sg13g2_fill_2
X_5074_ net399 VGND VPWR _0498_ videogen.test_lut_thingy.pixel_feeder_inst.row\[11\]\[1\]
+ _0155_ sg13g2_dfrbpq_1
XFILLER_38_853 VPWR VGND sg13g2_fill_2
X_4025_ _1693_ _1644_ _1692_ _0661_ videogen.test_lut_thingy.gol_counter_reg\[0\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_374 VPWR VGND sg13g2_decap_8
XFILLER_37_363 VPWR VGND sg13g2_decap_8
XFILLER_37_396 VPWR VGND sg13g2_fill_2
XFILLER_12_208 VPWR VGND sg13g2_decap_8
XFILLER_40_539 VPWR VGND sg13g2_decap_8
X_4927_ net368 VGND VPWR _0355_ videogen.fancy_shader.n646\[9\] net634 sg13g2_dfrbpq_2
X_4858_ net123 VGND VPWR _0286_ videogen.test_lut_thingy.pixel_feeder_inst.row\[6\]\[3\]
+ _0017_ sg13g2_dfrbpq_1
X_3809_ _1474_ _1475_ _1476_ _1477_ _1478_ VPWR VGND sg13g2_nor4_1
XFILLER_21_797 VPWR VGND sg13g2_fill_1
X_4789_ net690 net743 _0219_ VPWR VGND sg13g2_nor2_1
Xheichips25_bagel_23 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_48_606 VPWR VGND sg13g2_fill_1
XFILLER_29_820 VPWR VGND sg13g2_decap_4
X_5044__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_43_300 VPWR VGND sg13g2_decap_8
XFILLER_28_396 VPWR VGND sg13g2_decap_8
XFILLER_12_731 VPWR VGND sg13g2_decap_4
XFILLER_34_62 VPWR VGND sg13g2_decap_4
XFILLER_15_1017 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_8_768 VPWR VGND sg13g2_fill_2
XFILLER_7_289 VPWR VGND sg13g2_decap_8
XFILLER_4_974 VPWR VGND sg13g2_decap_8
XFILLER_47_650 VPWR VGND sg13g2_decap_4
XFILLER_47_683 VPWR VGND sg13g2_fill_2
XFILLER_35_823 VPWR VGND sg13g2_fill_1
X_5097__302 VPWR VGND net302 sg13g2_tiehi
XFILLER_35_845 VPWR VGND sg13g2_decap_8
XFILLER_15_580 VPWR VGND sg13g2_decap_8
X_2973_ net775 videogen.test_lut_thingy.pixel_feeder_inst.row\[0\]\[1\] _0795_ _0310_
+ VPWR VGND sg13g2_mux2_1
X_4712_ net678 net732 _0142_ VPWR VGND sg13g2_nor2_1
X_4643_ net666 net718 _0073_ VPWR VGND sg13g2_nor2_1
XFILLER_30_594 VPWR VGND sg13g2_decap_4
X_4574_ net572 _2201_ _0627_ VPWR VGND sg13g2_nor2_1
X_3525_ _1194_ _1016_ _1192_ VPWR VGND sg13g2_nand2b_1
X_3456_ _1125_ net609 videogen.fancy_shader.video_x\[8\] VPWR VGND sg13g2_xnor2_1
X_3387_ videogen.fancy_shader.video_x\[6\] videogen.fancy_shader.video_x\[5\] videogen.fancy_shader.video_x\[7\]
+ _1057_ VPWR VGND _0926_ sg13g2_nand4_1
X_5126_ net185 VGND VPWR _0550_ videogen.test_lut_thingy.pixel_feeder_inst.row\[28\]\[0\]
+ _0198_ sg13g2_dfrbpq_1
X_5057_ net80 VGND VPWR _0485_ videogen.test_lut_thingy.pixel_feeder_inst.row\[38\]\[0\]
+ _0142_ sg13g2_dfrbpq_1
X_4008_ videogen.test_lut_thingy.pixel_feeder_inst.row\[47\]\[0\] net578 _1676_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_37_182 VPWR VGND sg13g2_fill_2
XFILLER_25_311 VPWR VGND sg13g2_fill_2
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_867 VPWR VGND sg13g2_decap_8
XFILLER_41_848 VPWR VGND sg13g2_fill_2
XFILLER_4_215 VPWR VGND sg13g2_decap_4
XFILLER_20_20 VPWR VGND sg13g2_fill_1
XFILLER_1_900 VPWR VGND sg13g2_decap_8
X_5144__45 VPWR VGND net45 sg13g2_tiehi
XFILLER_20_75 VPWR VGND sg13g2_fill_1
XFILLER_0_410 VPWR VGND sg13g2_fill_1
XFILLER_0_421 VPWR VGND sg13g2_decap_8
XFILLER_1_977 VPWR VGND sg13g2_decap_8
XFILLER_49_959 VPWR VGND sg13g2_decap_8
Xhold40 serialize.bit_cnt\[1\] VPWR VGND net445 sg13g2_dlygate4sd3_1
XFILLER_29_62 VPWR VGND sg13g2_decap_8
XFILLER_16_300 VPWR VGND sg13g2_decap_8
XFILLER_29_694 VPWR VGND sg13g2_decap_4
XFILLER_16_366 VPWR VGND sg13g2_fill_2
XFILLER_17_867 VPWR VGND sg13g2_decap_4
XFILLER_43_163 VPWR VGND sg13g2_fill_1
XFILLER_31_314 VPWR VGND sg13g2_fill_1
XFILLER_31_325 VPWR VGND sg13g2_decap_4
XFILLER_32_859 VPWR VGND sg13g2_fill_1
X_4992__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_8_543 VPWR VGND sg13g2_fill_1
XFILLER_12_583 VPWR VGND sg13g2_fill_2
X_3310_ videogen.fancy_shader.n646\[3\] videogen.fancy_shader.video_x\[3\] _1000_
+ VPWR VGND sg13g2_nor2_1
X_4290_ VPWR VGND _1940_ _1926_ _1938_ _1928_ _1952_ _1929_ sg13g2_a221oi_1
X_3241_ videogen.test_lut_thingy.pixel_feeder_inst.v_pix\[4\] _0950_ _0951_ VPWR VGND
+ sg13g2_nor2_1
X_4964__317 VPWR VGND net317 sg13g2_tiehi
X_3172_ _0900_ _0899_ _0901_ VPWR VGND sg13g2_nor2b_2
XFILLER_48_970 VPWR VGND sg13g2_decap_8
XFILLER_23_859 VPWR VGND sg13g2_fill_1
X_2956_ videogen.test_lut_thingy.pixel_feeder_inst.row\[19\]\[3\] net760 _0792_ _0345_
+ VPWR VGND sg13g2_mux2_1
X_2887_ net759 videogen.test_lut_thingy.pixel_feeder_inst.row\[50\]\[3\] _0775_ _0440_
+ VPWR VGND sg13g2_mux2_1
X_4626_ net663 net715 _0056_ VPWR VGND sg13g2_nor2_1
X_4557_ _2153_ _2169_ _2151_ _2186_ VPWR VGND sg13g2_nand3_1
X_4488_ _2121_ _2118_ _2120_ VPWR VGND sg13g2_xnor2_1
X_3508_ net544 _1176_ _1177_ VPWR VGND sg13g2_nor2_1
X_3439_ _1108_ videogen.fancy_shader.video_y\[9\] videogen.fancy_shader.n646\[9\]
+ VPWR VGND sg13g2_xnor2_1
X_5109_ net252 VGND VPWR _0533_ videogen.test_lut_thingy.pixel_feeder_inst.row\[33\]\[3\]
+ _0181_ sg13g2_dfrbpq_1
XFILLER_38_480 VPWR VGND sg13g2_decap_4
XFILLER_25_130 VPWR VGND sg13g2_fill_1
XFILLER_26_686 VPWR VGND sg13g2_fill_2
XFILLER_26_697 VPWR VGND sg13g2_fill_2
XFILLER_40_166 VPWR VGND sg13g2_fill_2
XFILLER_31_52 VPWR VGND sg13g2_decap_4
Xoutput6 net6 tmds_r VPWR VGND sg13g2_buf_1
XFILLER_5_557 VPWR VGND sg13g2_decap_8
XFILLER_31_96 VPWR VGND sg13g2_decap_8
XFILLER_1_774 VPWR VGND sg13g2_decap_8
XFILLER_0_295 VPWR VGND sg13g2_fill_1
XFILLER_37_929 VPWR VGND sg13g2_decap_4
XFILLER_36_417 VPWR VGND sg13g2_fill_2
XFILLER_36_428 VPWR VGND sg13g2_fill_2
X_5020__204 VPWR VGND net204 sg13g2_tiehi
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_44_494 VPWR VGND sg13g2_fill_2
X_3790_ videogen.test_lut_thingy.pixel_feeder_inst.row\[58\]\[1\] net554 _1459_ VPWR
+ VGND sg13g2_nor2_1
X_2810_ net752 videogen.test_lut_thingy.pixel_feeder_inst.row\[15\]\[3\] _0754_ _0496_
+ VPWR VGND sg13g2_mux2_1
X_2741_ _0733_ _0737_ _0738_ VPWR VGND sg13g2_nor2_2
XFILLER_8_362 VPWR VGND sg13g2_fill_2
XFILLER_9_896 VPWR VGND sg13g2_decap_8
X_2672_ _0714_ _0716_ _0717_ VPWR VGND sg13g2_nor2b_2
X_4411_ _2055_ _2051_ _0913_ _2040_ _2015_ VPWR VGND sg13g2_a22oi_1
X_4342_ VGND VPWR _0860_ _0864_ _1993_ _1992_ sg13g2_a21oi_1
X_4273_ _1933_ VPWR _1935_ VGND _1914_ _1923_ sg13g2_o21ai_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_3224_ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[3\] VPWR _0938_ VGND
+ videogen.test_lut_thingy.pixel_feeder_inst.v_counter\[0\] _0820_ sg13g2_o21ai_1
.ends

