module heichips25_bagel (clk,
    ena,
    rst_n,
    tmds_b,
    tmds_clk,
    tmds_g,
    tmds_r,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 output tmds_b;
 output tmds_clk;
 output tmds_g;
 output tmds_r;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire clk_regs;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire \blue_tmds_par[0] ;
 wire \blue_tmds_par[1] ;
 wire \blue_tmds_par[2] ;
 wire \blue_tmds_par[3] ;
 wire \blue_tmds_par[5] ;
 wire \blue_tmds_par[6] ;
 wire \blue_tmds_par[7] ;
 wire \blue_tmds_par[8] ;
 wire \blue_tmds_par[9] ;
 wire clk_video;
 wire \clockdiv.q0 ;
 wire \clockdiv.q1 ;
 wire \clockdiv.q2 ;
 wire \clockdiv.q2temp ;
 wire display_enable;
 wire \green_tmds_par[0] ;
 wire \green_tmds_par[1] ;
 wire \green_tmds_par[2] ;
 wire \green_tmds_par[6] ;
 wire \green_tmds_par[7] ;
 wire \green_tmds_par[8] ;
 wire \green_tmds_par[9] ;
 wire hsync;
 wire \red_tmds_par[0] ;
 wire \red_tmds_par[1] ;
 wire \red_tmds_par[2] ;
 wire \red_tmds_par[3] ;
 wire \red_tmds_par[4] ;
 wire \red_tmds_par[5] ;
 wire \red_tmds_par[6] ;
 wire \red_tmds_par[7] ;
 wire \red_tmds_par[8] ;
 wire \red_tmds_par[9] ;
 wire \serialize.bit_cnt[0] ;
 wire \serialize.bit_cnt[1] ;
 wire \serialize.n410 ;
 wire \serialize.n411[0] ;
 wire \serialize.n411[1] ;
 wire \serialize.n411[2] ;
 wire \serialize.n411[3] ;
 wire \serialize.n411[4] ;
 wire \serialize.n411[5] ;
 wire \serialize.n411[6] ;
 wire \serialize.n411[7] ;
 wire \serialize.n414[0] ;
 wire \serialize.n414[1] ;
 wire \serialize.n414[2] ;
 wire \serialize.n414[3] ;
 wire \serialize.n414[4] ;
 wire \serialize.n414[5] ;
 wire \serialize.n414[6] ;
 wire \serialize.n414[7] ;
 wire \serialize.n417[0] ;
 wire \serialize.n417[1] ;
 wire \serialize.n417[2] ;
 wire \serialize.n417[3] ;
 wire \serialize.n417[4] ;
 wire \serialize.n417[5] ;
 wire \serialize.n417[6] ;
 wire \serialize.n417[7] ;
 wire \serialize.n420[0] ;
 wire \serialize.n420[1] ;
 wire \serialize.n420[2] ;
 wire \serialize.n420[3] ;
 wire \serialize.n420[4] ;
 wire \serialize.n420[6] ;
 wire \serialize.n427[0] ;
 wire \serialize.n427[1] ;
 wire \serialize.n427[2] ;
 wire \serialize.n427[3] ;
 wire \serialize.n427[4] ;
 wire \serialize.n427[5] ;
 wire \serialize.n427[6] ;
 wire \serialize.n427[7] ;
 wire \serialize.n427[8] ;
 wire \serialize.n427[9] ;
 wire \serialize.n428[0] ;
 wire \serialize.n428[1] ;
 wire \serialize.n428[2] ;
 wire \serialize.n428[3] ;
 wire \serialize.n428[4] ;
 wire \serialize.n428[5] ;
 wire \serialize.n428[6] ;
 wire \serialize.n428[7] ;
 wire \serialize.n428[8] ;
 wire \serialize.n428[9] ;
 wire \serialize.n429[0] ;
 wire \serialize.n429[1] ;
 wire \serialize.n429[2] ;
 wire \serialize.n429[3] ;
 wire \serialize.n429[4] ;
 wire \serialize.n429[5] ;
 wire \serialize.n429[6] ;
 wire \serialize.n429[7] ;
 wire \serialize.n429[8] ;
 wire \serialize.n429[9] ;
 wire \serialize.n431[0] ;
 wire \serialize.n431[1] ;
 wire \serialize.n431[2] ;
 wire \serialize.n431[3] ;
 wire \serialize.n431[4] ;
 wire \serialize.n431[5] ;
 wire \serialize.n431[6] ;
 wire \serialize.n433[0] ;
 wire \serialize.n433[1] ;
 wire \serialize.n450 ;
 wire \serialize.n452 ;
 wire \serialize.n453 ;
 wire \serialize.n455 ;
 wire \serialize.n456 ;
 wire \serialize.n458 ;
 wire \serialize.n459 ;
 wire \serialize.n461 ;
 wire net3;
 wire \tmds_blue.dc_balancing_reg[0] ;
 wire \tmds_blue.dc_balancing_reg[1] ;
 wire \tmds_blue.dc_balancing_reg[2] ;
 wire \tmds_blue.dc_balancing_reg[3] ;
 wire \tmds_blue.dc_balancing_reg[4] ;
 wire \tmds_blue.n100 ;
 wire \tmds_blue.n126 ;
 wire \tmds_blue.n132 ;
 wire \tmds_blue.n193 ;
 wire \tmds_blue.vsync ;
 wire net4;
 wire net5;
 wire \tmds_green.dc_balancing_reg[0] ;
 wire \tmds_green.dc_balancing_reg[1] ;
 wire \tmds_green.dc_balancing_reg[2] ;
 wire \tmds_green.dc_balancing_reg[3] ;
 wire \tmds_green.dc_balancing_reg[4] ;
 wire \tmds_green.n100 ;
 wire \tmds_green.n126 ;
 wire \tmds_green.n132 ;
 wire net6;
 wire \tmds_red.dc_balancing_reg[0] ;
 wire \tmds_red.dc_balancing_reg[1] ;
 wire \tmds_red.dc_balancing_reg[2] ;
 wire \tmds_red.dc_balancing_reg[3] ;
 wire \tmds_red.dc_balancing_reg[4] ;
 wire \tmds_red.n100 ;
 wire \tmds_red.n102 ;
 wire \tmds_red.n114 ;
 wire \tmds_red.n126 ;
 wire \tmds_red.n132 ;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net7;
 wire net28;
 wire net8;
 wire net9;
 wire net10;
 wire net29;
 wire net30;
 wire net31;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \videogen.fancy_shader.n646[0] ;
 wire \videogen.fancy_shader.n646[1] ;
 wire \videogen.fancy_shader.n646[2] ;
 wire \videogen.fancy_shader.n646[3] ;
 wire \videogen.fancy_shader.n646[4] ;
 wire \videogen.fancy_shader.n646[5] ;
 wire \videogen.fancy_shader.n646[6] ;
 wire \videogen.fancy_shader.n646[7] ;
 wire \videogen.fancy_shader.n646[8] ;
 wire \videogen.fancy_shader.n646[9] ;
 wire \videogen.fancy_shader.video_x[0] ;
 wire \videogen.fancy_shader.video_x[1] ;
 wire \videogen.fancy_shader.video_x[2] ;
 wire \videogen.fancy_shader.video_x[3] ;
 wire \videogen.fancy_shader.video_x[4] ;
 wire \videogen.fancy_shader.video_x[5] ;
 wire \videogen.fancy_shader.video_x[6] ;
 wire \videogen.fancy_shader.video_x[7] ;
 wire \videogen.fancy_shader.video_x[8] ;
 wire \videogen.fancy_shader.video_x[9] ;
 wire \videogen.fancy_shader.video_y[0] ;
 wire \videogen.fancy_shader.video_y[1] ;
 wire \videogen.fancy_shader.video_y[2] ;
 wire \videogen.fancy_shader.video_y[3] ;
 wire \videogen.fancy_shader.video_y[4] ;
 wire \videogen.fancy_shader.video_y[5] ;
 wire \videogen.fancy_shader.video_y[6] ;
 wire \videogen.fancy_shader.video_y[7] ;
 wire \videogen.fancy_shader.video_y[8] ;
 wire \videogen.fancy_shader.video_y[9] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[0] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[1] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[2] ;
 wire \videogen.test_lut_thingy.gol_counter_reg[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.state[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ;
 wire \videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net1;
 wire net2;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;

 sg13g2_inv_1 _2576_ (.Y(_0632_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ));
 sg13g2_inv_1 _2577_ (.Y(_0633_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ));
 sg13g2_inv_1 _2578_ (.Y(_0634_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ));
 sg13g2_inv_1 _2579_ (.Y(_0635_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ));
 sg13g2_inv_1 _2580_ (.Y(_0636_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ));
 sg13g2_inv_1 _2581_ (.Y(_0637_),
    .A(\videogen.fancy_shader.video_y[9] ));
 sg13g2_inv_1 _2582_ (.Y(_0638_),
    .A(\videogen.fancy_shader.video_y[8] ));
 sg13g2_inv_1 _2583_ (.Y(_0639_),
    .A(\videogen.fancy_shader.video_y[7] ));
 sg13g2_inv_1 _2584_ (.Y(_0640_),
    .A(\videogen.fancy_shader.video_y[2] ));
 sg13g2_inv_1 _2585_ (.Y(_0641_),
    .A(\videogen.fancy_shader.n646[9] ));
 sg13g2_inv_2 _2586_ (.Y(_0642_),
    .A(\videogen.fancy_shader.n646[7] ));
 sg13g2_inv_1 _2587_ (.Y(_0643_),
    .A(\videogen.fancy_shader.n646[0] ));
 sg13g2_inv_1 _2588_ (.Y(_0644_),
    .A(net611));
 sg13g2_inv_4 _2589_ (.A(net614),
    .Y(_0645_));
 sg13g2_inv_2 _2590_ (.Y(_0646_),
    .A(net619));
 sg13g2_inv_2 _2591_ (.Y(_0647_),
    .A(net628));
 sg13g2_inv_1 _2592_ (.Y(_0648_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ));
 sg13g2_inv_1 _2593_ (.Y(_0649_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ));
 sg13g2_inv_1 _2594_ (.Y(_0650_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ));
 sg13g2_inv_2 _2595_ (.Y(_0651_),
    .A(net629));
 sg13g2_inv_1 _2596_ (.Y(_0652_),
    .A(\tmds_green.dc_balancing_reg[1] ));
 sg13g2_inv_1 _2597_ (.Y(_0653_),
    .A(\tmds_green.dc_balancing_reg[3] ));
 sg13g2_inv_4 _2598_ (.A(\tmds_green.dc_balancing_reg[4] ),
    .Y(_0654_));
 sg13g2_inv_1 _2599_ (.Y(_0655_),
    .A(\tmds_blue.dc_balancing_reg[4] ));
 sg13g2_inv_1 _2600_ (.Y(_0656_),
    .A(\tmds_blue.dc_balancing_reg[1] ));
 sg13g2_inv_1 _2601_ (.Y(_0657_),
    .A(\tmds_blue.dc_balancing_reg[3] ));
 sg13g2_inv_1 _2602_ (.Y(_0658_),
    .A(net796));
 sg13g2_inv_2 _2603_ (.Y(_0659_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ));
 sg13g2_inv_1 _2604_ (.Y(_0660_),
    .A(\videogen.test_lut_thingy.gol_counter_reg[1] ));
 sg13g2_inv_2 _2605_ (.Y(_0661_),
    .A(net2));
 sg13g2_inv_2 _2606_ (.Y(_0662_),
    .A(net1));
 sg13g2_inv_1 _2607_ (.Y(_0663_),
    .A(\tmds_red.n102 ));
 sg13g2_inv_1 _2608_ (.Y(_0664_),
    .A(\tmds_red.dc_balancing_reg[4] ));
 sg13g2_inv_1 _2609_ (.Y(_0665_),
    .A(\tmds_red.dc_balancing_reg[1] ));
 sg13g2_inv_1 _2610_ (.Y(_0666_),
    .A(\tmds_red.dc_balancing_reg[3] ));
 sg13g2_inv_1 _2611_ (.Y(_0667_),
    .A(hsync));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_inv_1 _2613_ (.Y(_0668_),
    .A(net414));
 sg13g2_inv_1 _2614_ (.Y(_0669_),
    .A(net417));
 sg13g2_inv_1 _2615_ (.Y(_0670_),
    .A(net418));
 sg13g2_nand2_1 _2616_ (.Y(_0671_),
    .A(\serialize.bit_cnt[1] ),
    .B(net412));
 sg13g2_xor2_1 _2617_ (.B(net412),
    .A(net445),
    .X(\serialize.n433[1] ));
 sg13g2_nand2_1 _2618_ (.Y(_0672_),
    .A(net415),
    .B(_0671_));
 sg13g2_o21ai_1 _2619_ (.B1(_0672_),
    .Y(_0262_),
    .A1(net415),
    .A2(\serialize.n433[1] ));
 sg13g2_nand3_1 _2620_ (.B(\videogen.fancy_shader.video_y[6] ),
    .C(\videogen.fancy_shader.video_y[5] ),
    .A(\videogen.fancy_shader.video_y[7] ),
    .Y(_0673_));
 sg13g2_nor3_1 _2621_ (.A(\videogen.fancy_shader.video_y[9] ),
    .B(_0638_),
    .C(_0673_),
    .Y(_0674_));
 sg13g2_nor2b_1 _2622_ (.A(\videogen.fancy_shader.video_y[4] ),
    .B_N(_0674_),
    .Y(_0675_));
 sg13g2_nor4_1 _2623_ (.A(\videogen.fancy_shader.video_y[3] ),
    .B(\videogen.fancy_shader.video_y[2] ),
    .C(\videogen.fancy_shader.video_y[1] ),
    .D(net608),
    .Y(_0676_));
 sg13g2_and2_1 _2624_ (.A(_0675_),
    .B(_0676_),
    .X(_0677_));
 sg13g2_nor3_1 _2625_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(\videogen.fancy_shader.video_x[5] ),
    .C(\videogen.fancy_shader.video_x[4] ),
    .Y(_0678_));
 sg13g2_nor3_1 _2626_ (.A(_0651_),
    .B(\videogen.fancy_shader.video_x[3] ),
    .C(\videogen.fancy_shader.video_x[2] ),
    .Y(_0679_));
 sg13g2_nor2b_2 _2627_ (.A(\videogen.fancy_shader.video_x[8] ),
    .B_N(\videogen.fancy_shader.video_x[9] ),
    .Y(_0680_));
 sg13g2_nor2_1 _2628_ (.A(\videogen.fancy_shader.video_x[1] ),
    .B(\videogen.fancy_shader.video_x[0] ),
    .Y(_0681_));
 sg13g2_nand4_1 _2629_ (.B(_0679_),
    .C(_0680_),
    .A(_0678_),
    .Y(_0682_),
    .D(_0681_));
 sg13g2_inv_2 _2630_ (.Y(_0683_),
    .A(_0682_));
 sg13g2_nor2_2 _2631_ (.A(_0677_),
    .B(_0682_),
    .Y(_0684_));
 sg13g2_nand2_2 _2632_ (.Y(_0685_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .B(_0684_));
 sg13g2_nor2_1 _2633_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .B(net628),
    .Y(_0686_));
 sg13g2_or2_1 _2634_ (.X(_0687_),
    .B(net628),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ));
 sg13g2_nor2_1 _2635_ (.A(net619),
    .B(net587),
    .Y(_0688_));
 sg13g2_nor3_1 _2636_ (.A(net614),
    .B(net620),
    .C(net585),
    .Y(_0689_));
 sg13g2_xnor2_1 _2637_ (.Y(_0690_),
    .A(net615),
    .B(_0688_));
 sg13g2_nand2_2 _2638_ (.Y(_0691_),
    .A(_0685_),
    .B(_0690_));
 sg13g2_and2_1 _2639_ (.A(_0644_),
    .B(_0689_),
    .X(_0692_));
 sg13g2_xnor2_1 _2640_ (.Y(_0693_),
    .A(net611),
    .B(_0689_));
 sg13g2_nand2b_2 _2641_ (.Y(_0694_),
    .B(_0692_),
    .A_N(net610));
 sg13g2_xnor2_1 _2642_ (.Y(_0695_),
    .A(net610),
    .B(_0692_));
 sg13g2_nand2_1 _2643_ (.Y(_0696_),
    .A(_0685_),
    .B(_0695_));
 sg13g2_nand2_1 _2644_ (.Y(_0697_),
    .A(_0685_),
    .B(_0693_));
 sg13g2_nand3_1 _2645_ (.B(_0693_),
    .C(_0695_),
    .A(_0685_),
    .Y(_0698_));
 sg13g2_nor2b_2 _2646_ (.A(_0698_),
    .B_N(net545),
    .Y(_0699_));
 sg13g2_nand2b_2 _2647_ (.Y(_0700_),
    .B(net545),
    .A_N(_0698_));
 sg13g2_and2_1 _2648_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .B(net628),
    .X(_0701_));
 sg13g2_nand2_2 _2649_ (.Y(_0702_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .B(net628));
 sg13g2_nor2_1 _2650_ (.A(net593),
    .B(net583),
    .Y(_0703_));
 sg13g2_and2_1 _2651_ (.A(_0685_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nand2_1 _2652_ (.Y(_0705_),
    .A(_0685_),
    .B(_0703_));
 sg13g2_nor3_1 _2653_ (.A(_0647_),
    .B(net595),
    .C(_0684_),
    .Y(_0706_));
 sg13g2_nand3_1 _2654_ (.B(_0705_),
    .C(_0706_),
    .A(net619),
    .Y(_0707_));
 sg13g2_nor2_2 _2655_ (.A(_0700_),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_mux2_1 _2656_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .A1(net753),
    .S(_0708_),
    .X(_0631_));
 sg13g2_mux2_1 _2657_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .A1(net763),
    .S(_0708_),
    .X(_0630_));
 sg13g2_mux2_1 _2658_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .A1(net773),
    .S(_0708_),
    .X(_0629_));
 sg13g2_mux2_1 _2659_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .A1(net784),
    .S(_0708_),
    .X(_0628_));
 sg13g2_xnor2_1 _2660_ (.Y(_0709_),
    .A(net619),
    .B(net593));
 sg13g2_nand3b_1 _2661_ (.B(_0709_),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .Y(_0710_),
    .A_N(_0684_));
 sg13g2_nor2_2 _2662_ (.A(net573),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_or2_1 _2663_ (.X(_0712_),
    .B(_0710_),
    .A(net573));
 sg13g2_nand2_2 _2664_ (.Y(_0713_),
    .A(_0699_),
    .B(_0711_));
 sg13g2_mux2_1 _2665_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .S(_0713_),
    .X(_0609_));
 sg13g2_mux2_1 _2666_ (.A0(net763),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .S(_0713_),
    .X(_0608_));
 sg13g2_mux2_1 _2667_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .S(_0713_),
    .X(_0607_));
 sg13g2_mux2_1 _2668_ (.A0(net785),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .S(_0713_),
    .X(_0606_));
 sg13g2_or2_1 _2669_ (.X(_0714_),
    .B(_0698_),
    .A(net545));
 sg13g2_nand2_1 _2670_ (.Y(_0715_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .B(_0688_));
 sg13g2_nand2_2 _2671_ (.Y(_0716_),
    .A(_0685_),
    .B(_0715_));
 sg13g2_nor2b_2 _2672_ (.A(_0714_),
    .B_N(_0716_),
    .Y(_0717_));
 sg13g2_mux2_1 _2673_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .A1(net753),
    .S(_0717_),
    .X(_0605_));
 sg13g2_mux2_1 _2674_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .A1(net762),
    .S(_0717_),
    .X(_0604_));
 sg13g2_mux2_1 _2675_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .A1(net773),
    .S(_0717_),
    .X(_0603_));
 sg13g2_mux2_1 _2676_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .A1(net784),
    .S(_0717_),
    .X(_0602_));
 sg13g2_nor2_2 _2677_ (.A(_0693_),
    .B(_0696_),
    .Y(_0718_));
 sg13g2_nand2b_2 _2678_ (.Y(_0719_),
    .B(_0718_),
    .A_N(net545));
 sg13g2_and3_2 _2679_ (.X(_0720_),
    .A(_0646_),
    .B(_0704_),
    .C(_0706_));
 sg13g2_nand2b_2 _2680_ (.Y(_0721_),
    .B(_0720_),
    .A_N(_0719_));
 sg13g2_mux2_1 _2681_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ),
    .S(_0721_),
    .X(_0601_));
 sg13g2_mux2_1 _2682_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .S(_0721_),
    .X(_0600_));
 sg13g2_mux2_1 _2683_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ),
    .S(_0721_),
    .X(_0599_));
 sg13g2_mux2_1 _2684_ (.A0(net792),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ),
    .S(_0721_),
    .X(_0598_));
 sg13g2_nor4_2 _2685_ (.A(net619),
    .B(net628),
    .C(net595),
    .Y(_0722_),
    .D(_0705_));
 sg13g2_nand2b_2 _2686_ (.Y(_0723_),
    .B(_0722_),
    .A_N(_0719_));
 sg13g2_mux2_1 _2687_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .S(_0723_),
    .X(_0597_));
 sg13g2_mux2_1 _2688_ (.A0(net770),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .S(_0723_),
    .X(_0596_));
 sg13g2_mux2_1 _2689_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .S(_0723_),
    .X(_0595_));
 sg13g2_mux2_1 _2690_ (.A0(net792),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .S(_0723_),
    .X(_0594_));
 sg13g2_nor2_2 _2691_ (.A(_0712_),
    .B(_0719_),
    .Y(_0724_));
 sg13g2_mux2_1 _2692_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .A1(net760),
    .S(_0724_),
    .X(_0593_));
 sg13g2_mux2_1 _2693_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .A1(net770),
    .S(_0724_),
    .X(_0592_));
 sg13g2_mux2_1 _2694_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .A1(net782),
    .S(_0724_),
    .X(_0591_));
 sg13g2_mux2_1 _2695_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .A1(net793),
    .S(_0724_),
    .X(_0590_));
 sg13g2_nor2b_2 _2696_ (.A(_0714_),
    .B_N(_0722_),
    .Y(_0725_));
 sg13g2_mux2_1 _2697_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .A1(net754),
    .S(_0725_),
    .X(_0589_));
 sg13g2_mux2_1 _2698_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .A1(net762),
    .S(_0725_),
    .X(_0588_));
 sg13g2_mux2_1 _2699_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .A1(net775),
    .S(_0725_),
    .X(_0587_));
 sg13g2_mux2_1 _2700_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .A1(net786),
    .S(_0725_),
    .X(_0586_));
 sg13g2_nand3_1 _2701_ (.B(_0704_),
    .C(_0706_),
    .A(net619),
    .Y(_0726_));
 sg13g2_nor2_2 _2702_ (.A(_0719_),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_mux2_1 _2703_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .A1(net760),
    .S(_0727_),
    .X(_0585_));
 sg13g2_mux2_1 _2704_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .A1(net770),
    .S(_0727_),
    .X(_0584_));
 sg13g2_mux2_1 _2705_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .A1(net782),
    .S(_0727_),
    .X(_0583_));
 sg13g2_mux2_1 _2706_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .A1(net792),
    .S(_0727_),
    .X(_0582_));
 sg13g2_nand4_1 _2707_ (.B(_0647_),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .A(net619),
    .Y(_0728_),
    .D(_0704_));
 sg13g2_nor2_2 _2708_ (.A(_0719_),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_mux2_1 _2709_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .A1(net760),
    .S(_0729_),
    .X(_0581_));
 sg13g2_mux2_1 _2710_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .A1(net770),
    .S(_0729_),
    .X(_0580_));
 sg13g2_mux2_1 _2711_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .A1(net782),
    .S(_0729_),
    .X(_0579_));
 sg13g2_mux2_1 _2712_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .A1(net792),
    .S(_0729_),
    .X(_0578_));
 sg13g2_nor2_2 _2713_ (.A(_0707_),
    .B(_0719_),
    .Y(_0730_));
 sg13g2_mux2_1 _2714_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .A1(net759),
    .S(_0730_),
    .X(_0577_));
 sg13g2_mux2_1 _2715_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .A1(net770),
    .S(_0730_),
    .X(_0576_));
 sg13g2_mux2_1 _2716_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .A1(net782),
    .S(_0730_),
    .X(_0575_));
 sg13g2_mux2_1 _2717_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .A1(net792),
    .S(_0730_),
    .X(_0574_));
 sg13g2_nand2b_2 _2718_ (.Y(_0731_),
    .B(_0716_),
    .A_N(_0719_));
 sg13g2_mux2_1 _2719_ (.A0(net760),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .S(_0731_),
    .X(_0573_));
 sg13g2_mux2_1 _2720_ (.A0(net772),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .S(_0731_),
    .X(_0572_));
 sg13g2_mux2_1 _2721_ (.A0(net782),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .S(_0731_),
    .X(_0571_));
 sg13g2_mux2_1 _2722_ (.A0(net792),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .S(_0731_),
    .X(_0570_));
 sg13g2_and2_1 _2723_ (.A(net546),
    .B(_0718_),
    .X(_0732_));
 sg13g2_nand2_2 _2724_ (.Y(_0733_),
    .A(net546),
    .B(_0718_));
 sg13g2_nand2_2 _2725_ (.Y(_0734_),
    .A(_0720_),
    .B(_0732_));
 sg13g2_mux2_1 _2726_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .S(_0734_),
    .X(_0569_));
 sg13g2_mux2_1 _2727_ (.A0(net762),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .S(_0734_),
    .X(_0568_));
 sg13g2_mux2_1 _2728_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .S(_0734_),
    .X(_0567_));
 sg13g2_mux2_1 _2729_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ),
    .S(_0734_),
    .X(_0566_));
 sg13g2_nand2_2 _2730_ (.Y(_0735_),
    .A(_0722_),
    .B(_0732_));
 sg13g2_mux2_1 _2731_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .S(_0735_),
    .X(_0565_));
 sg13g2_mux2_1 _2732_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .S(_0735_),
    .X(_0564_));
 sg13g2_mux2_1 _2733_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .S(_0735_),
    .X(_0563_));
 sg13g2_mux2_1 _2734_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .S(_0735_),
    .X(_0562_));
 sg13g2_nand2_2 _2735_ (.Y(_0736_),
    .A(_0711_),
    .B(_0732_));
 sg13g2_mux2_1 _2736_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .S(_0736_),
    .X(_0561_));
 sg13g2_mux2_1 _2737_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .S(_0736_),
    .X(_0560_));
 sg13g2_mux2_1 _2738_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .S(_0736_),
    .X(_0559_));
 sg13g2_mux2_1 _2739_ (.A0(net794),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ),
    .S(_0736_),
    .X(_0558_));
 sg13g2_or2_1 _2740_ (.X(_0737_),
    .B(_0710_),
    .A(net585));
 sg13g2_nor2_2 _2741_ (.A(_0733_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_mux2_1 _2742_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ),
    .A1(net752),
    .S(_0738_),
    .X(_0557_));
 sg13g2_mux2_1 _2743_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .A1(net769),
    .S(_0738_),
    .X(_0556_));
 sg13g2_mux2_1 _2744_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ),
    .A1(net777),
    .S(_0738_),
    .X(_0555_));
 sg13g2_mux2_1 _2745_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .A1(net785),
    .S(_0738_),
    .X(_0554_));
 sg13g2_nor2_2 _2746_ (.A(_0726_),
    .B(_0733_),
    .Y(_0739_));
 sg13g2_mux2_1 _2747_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .A1(net759),
    .S(_0739_),
    .X(_0553_));
 sg13g2_mux2_1 _2748_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .A1(net770),
    .S(_0739_),
    .X(_0552_));
 sg13g2_mux2_1 _2749_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .A1(net781),
    .S(_0739_),
    .X(_0551_));
 sg13g2_mux2_1 _2750_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .A1(net791),
    .S(_0739_),
    .X(_0550_));
 sg13g2_nor2_2 _2751_ (.A(_0712_),
    .B(_0714_),
    .Y(_0740_));
 sg13g2_mux2_1 _2752_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .A1(net756),
    .S(_0740_),
    .X(_0549_));
 sg13g2_mux2_1 _2753_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .A1(net765),
    .S(_0740_),
    .X(_0548_));
 sg13g2_mux2_1 _2754_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .A1(net775),
    .S(_0740_),
    .X(_0547_));
 sg13g2_mux2_1 _2755_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .A1(net786),
    .S(_0740_),
    .X(_0546_));
 sg13g2_nor2_2 _2756_ (.A(_0707_),
    .B(_0733_),
    .Y(_0741_));
 sg13g2_mux2_1 _2757_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .A1(net756),
    .S(_0741_),
    .X(_0545_));
 sg13g2_mux2_1 _2758_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .A1(net771),
    .S(_0741_),
    .X(_0544_));
 sg13g2_mux2_1 _2759_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .A1(net777),
    .S(_0741_),
    .X(_0543_));
 sg13g2_mux2_1 _2760_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ),
    .A1(net788),
    .S(_0741_),
    .X(_0542_));
 sg13g2_nand2_2 _2761_ (.Y(_0742_),
    .A(_0716_),
    .B(_0732_));
 sg13g2_mux2_1 _2762_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .S(_0742_),
    .X(_0541_));
 sg13g2_mux2_1 _2763_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .S(_0742_),
    .X(_0540_));
 sg13g2_mux2_1 _2764_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .S(_0742_),
    .X(_0539_));
 sg13g2_mux2_1 _2765_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ),
    .S(_0742_),
    .X(_0538_));
 sg13g2_nor2_2 _2766_ (.A(_0695_),
    .B(_0697_),
    .Y(_0743_));
 sg13g2_nor3_2 _2767_ (.A(net545),
    .B(_0695_),
    .C(_0697_),
    .Y(_0744_));
 sg13g2_nand2b_2 _2768_ (.Y(_0745_),
    .B(_0743_),
    .A_N(net545));
 sg13g2_nand2_2 _2769_ (.Y(_0746_),
    .A(_0720_),
    .B(_0744_));
 sg13g2_mux2_1 _2770_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .S(_0746_),
    .X(_0537_));
 sg13g2_mux2_1 _2771_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .S(_0746_),
    .X(_0536_));
 sg13g2_mux2_1 _2772_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .S(_0746_),
    .X(_0535_));
 sg13g2_mux2_1 _2773_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .S(_0746_),
    .X(_0534_));
 sg13g2_nand2_2 _2774_ (.Y(_0747_),
    .A(_0722_),
    .B(_0744_));
 sg13g2_mux2_1 _2775_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .S(_0747_),
    .X(_0533_));
 sg13g2_mux2_1 _2776_ (.A0(net767),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .S(_0747_),
    .X(_0532_));
 sg13g2_mux2_1 _2777_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .S(_0747_),
    .X(_0531_));
 sg13g2_mux2_1 _2778_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .S(_0747_),
    .X(_0530_));
 sg13g2_nor2_2 _2779_ (.A(_0712_),
    .B(_0745_),
    .Y(_0748_));
 sg13g2_mux2_1 _2780_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .A1(net757),
    .S(_0748_),
    .X(_0529_));
 sg13g2_mux2_1 _2781_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .A1(net767),
    .S(_0748_),
    .X(_0528_));
 sg13g2_mux2_1 _2782_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .A1(net779),
    .S(_0748_),
    .X(_0527_));
 sg13g2_mux2_1 _2783_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .A1(net790),
    .S(_0748_),
    .X(_0526_));
 sg13g2_nor2_2 _2784_ (.A(_0737_),
    .B(_0745_),
    .Y(_0749_));
 sg13g2_mux2_1 _2785_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .A1(net752),
    .S(_0749_),
    .X(_0525_));
 sg13g2_mux2_1 _2786_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .A1(net767),
    .S(_0749_),
    .X(_0524_));
 sg13g2_mux2_1 _2787_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ),
    .A1(net774),
    .S(_0749_),
    .X(_0523_));
 sg13g2_mux2_1 _2788_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ),
    .A1(net785),
    .S(_0749_),
    .X(_0522_));
 sg13g2_nor2_2 _2789_ (.A(_0726_),
    .B(_0745_),
    .Y(_0750_));
 sg13g2_mux2_1 _2790_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .A1(net758),
    .S(_0750_),
    .X(_0521_));
 sg13g2_mux2_1 _2791_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .A1(net768),
    .S(_0750_),
    .X(_0520_));
 sg13g2_mux2_1 _2792_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .A1(net779),
    .S(_0750_),
    .X(_0519_));
 sg13g2_mux2_1 _2793_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .A1(net789),
    .S(_0750_),
    .X(_0518_));
 sg13g2_nor2_2 _2794_ (.A(_0728_),
    .B(_0745_),
    .Y(_0751_));
 sg13g2_mux2_1 _2795_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .A1(net758),
    .S(_0751_),
    .X(_0517_));
 sg13g2_mux2_1 _2796_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .A1(net768),
    .S(_0751_),
    .X(_0516_));
 sg13g2_mux2_1 _2797_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .A1(net780),
    .S(_0751_),
    .X(_0515_));
 sg13g2_mux2_1 _2798_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .A1(net789),
    .S(_0751_),
    .X(_0514_));
 sg13g2_nor2_2 _2799_ (.A(_0700_),
    .B(_0728_),
    .Y(_0752_));
 sg13g2_mux2_1 _2800_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .A1(net753),
    .S(_0752_),
    .X(_0504_));
 sg13g2_mux2_1 _2801_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .A1(net762),
    .S(_0752_),
    .X(_0503_));
 sg13g2_mux2_1 _2802_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .A1(net773),
    .S(_0752_),
    .X(_0502_));
 sg13g2_mux2_1 _2803_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .A1(net784),
    .S(_0752_),
    .X(_0501_));
 sg13g2_nor2_2 _2804_ (.A(_0700_),
    .B(_0737_),
    .Y(_0753_));
 sg13g2_mux2_1 _2805_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .A1(net753),
    .S(_0753_),
    .X(_0500_));
 sg13g2_mux2_1 _2806_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .A1(net762),
    .S(_0753_),
    .X(_0499_));
 sg13g2_mux2_1 _2807_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ),
    .A1(net773),
    .S(_0753_),
    .X(_0498_));
 sg13g2_mux2_1 _2808_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .A1(net784),
    .S(_0753_),
    .X(_0497_));
 sg13g2_nand2_2 _2809_ (.Y(_0754_),
    .A(_0699_),
    .B(_0716_));
 sg13g2_mux2_1 _2810_ (.A0(net752),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .S(_0754_),
    .X(_0496_));
 sg13g2_mux2_1 _2811_ (.A0(net763),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .S(_0754_),
    .X(_0495_));
 sg13g2_mux2_1 _2812_ (.A0(net774),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .S(_0754_),
    .X(_0494_));
 sg13g2_mux2_1 _2813_ (.A0(net785),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .S(_0754_),
    .X(_0493_));
 sg13g2_nor2_2 _2814_ (.A(_0714_),
    .B(_0737_),
    .Y(_0755_));
 sg13g2_mux2_1 _2815_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ),
    .A1(net754),
    .S(_0755_),
    .X(_0492_));
 sg13g2_mux2_1 _2816_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .A1(net765),
    .S(_0755_),
    .X(_0491_));
 sg13g2_mux2_1 _2817_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .A1(net775),
    .S(_0755_),
    .X(_0490_));
 sg13g2_mux2_1 _2818_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .A1(net786),
    .S(_0755_),
    .X(_0489_));
 sg13g2_nor2_2 _2819_ (.A(_0707_),
    .B(_0745_),
    .Y(_0756_));
 sg13g2_mux2_1 _2820_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .A1(net758),
    .S(_0756_),
    .X(_0488_));
 sg13g2_mux2_1 _2821_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .A1(net768),
    .S(_0756_),
    .X(_0487_));
 sg13g2_mux2_1 _2822_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .A1(net780),
    .S(_0756_),
    .X(_0486_));
 sg13g2_mux2_1 _2823_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .A1(net789),
    .S(_0756_),
    .X(_0485_));
 sg13g2_and2_1 _2824_ (.A(net545),
    .B(_0743_),
    .X(_0757_));
 sg13g2_nand2_2 _2825_ (.Y(_0758_),
    .A(net545),
    .B(_0743_));
 sg13g2_nand2_2 _2826_ (.Y(_0759_),
    .A(_0720_),
    .B(_0757_));
 sg13g2_mux2_1 _2827_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .S(_0759_),
    .X(_0484_));
 sg13g2_mux2_1 _2828_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .S(_0759_),
    .X(_0483_));
 sg13g2_mux2_1 _2829_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .S(_0759_),
    .X(_0482_));
 sg13g2_mux2_1 _2830_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .S(_0759_),
    .X(_0481_));
 sg13g2_nand2_2 _2831_ (.Y(_0760_),
    .A(_0699_),
    .B(_0720_));
 sg13g2_mux2_1 _2832_ (.A0(net753),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ),
    .S(_0760_),
    .X(_0480_));
 sg13g2_mux2_1 _2833_ (.A0(net762),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .S(_0760_),
    .X(_0479_));
 sg13g2_mux2_1 _2834_ (.A0(net773),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .S(_0760_),
    .X(_0478_));
 sg13g2_mux2_1 _2835_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ),
    .S(_0760_),
    .X(_0477_));
 sg13g2_nand2_2 _2836_ (.Y(_0761_),
    .A(_0722_),
    .B(_0757_));
 sg13g2_mux2_1 _2837_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .S(_0761_),
    .X(_0476_));
 sg13g2_mux2_1 _2838_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .S(_0761_),
    .X(_0475_));
 sg13g2_mux2_1 _2839_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ),
    .S(_0761_),
    .X(_0474_));
 sg13g2_mux2_1 _2840_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ),
    .S(_0761_),
    .X(_0473_));
 sg13g2_nand2_2 _2841_ (.Y(_0762_),
    .A(_0711_),
    .B(_0757_));
 sg13g2_mux2_1 _2842_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .S(_0762_),
    .X(_0472_));
 sg13g2_mux2_1 _2843_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .S(_0762_),
    .X(_0471_));
 sg13g2_mux2_1 _2844_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .S(_0762_),
    .X(_0470_));
 sg13g2_mux2_1 _2845_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .S(_0762_),
    .X(_0469_));
 sg13g2_nor2_2 _2846_ (.A(_0737_),
    .B(_0758_),
    .Y(_0763_));
 sg13g2_mux2_1 _2847_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .A1(net758),
    .S(_0763_),
    .X(_0468_));
 sg13g2_mux2_1 _2848_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .A1(net768),
    .S(_0763_),
    .X(_0467_));
 sg13g2_mux2_1 _2849_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .A1(net780),
    .S(_0763_),
    .X(_0466_));
 sg13g2_mux2_1 _2850_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .A1(net789),
    .S(_0763_),
    .X(_0465_));
 sg13g2_nor2_2 _2851_ (.A(_0726_),
    .B(_0758_),
    .Y(_0764_));
 sg13g2_nand2_1 _2852_ (.Y(_0765_),
    .A(net757),
    .B(_0764_));
 sg13g2_o21ai_1 _2853_ (.B1(_0765_),
    .Y(_0464_),
    .A1(_0632_),
    .A2(_0764_));
 sg13g2_mux2_1 _2854_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .A1(net767),
    .S(_0764_),
    .X(_0463_));
 sg13g2_mux2_1 _2855_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .A1(net779),
    .S(_0764_),
    .X(_0462_));
 sg13g2_mux2_1 _2856_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .A1(net790),
    .S(_0764_),
    .X(_0461_));
 sg13g2_nand2b_2 _2857_ (.Y(_0766_),
    .B(_0757_),
    .A_N(_0728_));
 sg13g2_mux2_1 _2858_ (.A0(net757),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .S(_0766_),
    .X(_0460_));
 sg13g2_mux2_1 _2859_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .S(_0766_),
    .X(_0459_));
 sg13g2_mux2_1 _2860_ (.A0(net780),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .S(_0766_),
    .X(_0458_));
 sg13g2_mux2_1 _2861_ (.A0(net790),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ),
    .S(_0766_),
    .X(_0457_));
 sg13g2_nor2_2 _2862_ (.A(_0707_),
    .B(_0758_),
    .Y(_0767_));
 sg13g2_mux2_1 _2863_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .A1(net757),
    .S(_0767_),
    .X(_0456_));
 sg13g2_mux2_1 _2864_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .A1(net767),
    .S(_0767_),
    .X(_0455_));
 sg13g2_mux2_1 _2865_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .A1(net779),
    .S(_0767_),
    .X(_0454_));
 sg13g2_mux2_1 _2866_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ),
    .A1(net790),
    .S(_0767_),
    .X(_0453_));
 sg13g2_nand2_2 _2867_ (.Y(_0768_),
    .A(_0716_),
    .B(_0757_));
 sg13g2_nor2_1 _2868_ (.A(net757),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_a21oi_1 _2869_ (.A1(_0633_),
    .A2(_0768_),
    .Y(_0452_),
    .B1(_0769_));
 sg13g2_mux2_1 _2870_ (.A0(net769),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .S(_0768_),
    .X(_0451_));
 sg13g2_mux2_1 _2871_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .S(_0768_),
    .X(_0450_));
 sg13g2_mux2_1 _2872_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .S(_0768_),
    .X(_0449_));
 sg13g2_o21ai_1 _2873_ (.B1(_0685_),
    .Y(_0770_),
    .A1(_0693_),
    .A2(_0695_));
 sg13g2_nor2b_2 _2874_ (.A(net546),
    .B_N(_0770_),
    .Y(_0771_));
 sg13g2_nand2b_2 _2875_ (.Y(_0772_),
    .B(_0770_),
    .A_N(net546));
 sg13g2_nand2_2 _2876_ (.Y(_0773_),
    .A(_0720_),
    .B(_0771_));
 sg13g2_mux2_1 _2877_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .S(_0773_),
    .X(_0448_));
 sg13g2_mux2_1 _2878_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .S(_0773_),
    .X(_0447_));
 sg13g2_mux2_1 _2879_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .S(_0773_),
    .X(_0446_));
 sg13g2_mux2_1 _2880_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .S(_0773_),
    .X(_0445_));
 sg13g2_nor2_2 _2881_ (.A(_0714_),
    .B(_0726_),
    .Y(_0774_));
 sg13g2_mux2_1 _2882_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .A1(net753),
    .S(_0774_),
    .X(_0444_));
 sg13g2_mux2_1 _2883_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .A1(net763),
    .S(_0774_),
    .X(_0443_));
 sg13g2_mux2_1 _2884_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .A1(net773),
    .S(_0774_),
    .X(_0442_));
 sg13g2_mux2_1 _2885_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .A1(net784),
    .S(_0774_),
    .X(_0441_));
 sg13g2_nand2_2 _2886_ (.Y(_0775_),
    .A(_0711_),
    .B(_0771_));
 sg13g2_mux2_1 _2887_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .S(_0775_),
    .X(_0440_));
 sg13g2_mux2_1 _2888_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .S(_0775_),
    .X(_0439_));
 sg13g2_mux2_1 _2889_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .S(_0775_),
    .X(_0438_));
 sg13g2_mux2_1 _2890_ (.A0(net792),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .S(_0775_),
    .X(_0437_));
 sg13g2_nor2_2 _2891_ (.A(_0737_),
    .B(_0772_),
    .Y(_0776_));
 sg13g2_mux2_1 _2892_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .A1(net759),
    .S(_0776_),
    .X(_0436_));
 sg13g2_mux2_1 _2893_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .A1(net771),
    .S(_0776_),
    .X(_0435_));
 sg13g2_mux2_1 _2894_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ),
    .A1(net781),
    .S(_0776_),
    .X(_0434_));
 sg13g2_mux2_1 _2895_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .A1(net791),
    .S(_0776_),
    .X(_0433_));
 sg13g2_nor2_2 _2896_ (.A(_0726_),
    .B(_0772_),
    .Y(_0777_));
 sg13g2_mux2_1 _2897_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .A1(net755),
    .S(_0777_),
    .X(_0432_));
 sg13g2_mux2_1 _2898_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .A1(net764),
    .S(_0777_),
    .X(_0431_));
 sg13g2_mux2_1 _2899_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .A1(net777),
    .S(_0777_),
    .X(_0430_));
 sg13g2_mux2_1 _2900_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ),
    .A1(net788),
    .S(_0777_),
    .X(_0429_));
 sg13g2_nor2_2 _2901_ (.A(_0728_),
    .B(_0772_),
    .Y(_0778_));
 sg13g2_mux2_1 _2902_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .A1(net755),
    .S(_0778_),
    .X(_0428_));
 sg13g2_mux2_1 _2903_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .A1(net765),
    .S(_0778_),
    .X(_0427_));
 sg13g2_mux2_1 _2904_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .A1(net777),
    .S(_0778_),
    .X(_0426_));
 sg13g2_mux2_1 _2905_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .A1(net788),
    .S(_0778_),
    .X(_0425_));
 sg13g2_nor2_2 _2906_ (.A(_0707_),
    .B(_0772_),
    .Y(_0779_));
 sg13g2_mux2_1 _2907_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .A1(net755),
    .S(_0779_),
    .X(_0424_));
 sg13g2_mux2_1 _2908_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .A1(net765),
    .S(_0779_),
    .X(_0423_));
 sg13g2_mux2_1 _2909_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .A1(net778),
    .S(_0779_),
    .X(_0422_));
 sg13g2_mux2_1 _2910_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .A1(net788),
    .S(_0779_),
    .X(_0421_));
 sg13g2_nand2_2 _2911_ (.Y(_0780_),
    .A(_0716_),
    .B(_0771_));
 sg13g2_mux2_1 _2912_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .S(_0780_),
    .X(_0420_));
 sg13g2_mux2_1 _2913_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .S(_0780_),
    .X(_0419_));
 sg13g2_mux2_1 _2914_ (.A0(net777),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .S(_0780_),
    .X(_0418_));
 sg13g2_mux2_1 _2915_ (.A0(net788),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ),
    .S(_0780_),
    .X(_0417_));
 sg13g2_and2_1 _2916_ (.A(net546),
    .B(_0770_),
    .X(_0781_));
 sg13g2_nand2_2 _2917_ (.Y(_0782_),
    .A(_0720_),
    .B(_0781_));
 sg13g2_mux2_1 _2918_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .S(_0782_),
    .X(_0416_));
 sg13g2_mux2_1 _2919_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .S(_0782_),
    .X(_0415_));
 sg13g2_mux2_1 _2920_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .S(_0782_),
    .X(_0414_));
 sg13g2_mux2_1 _2921_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ),
    .S(_0782_),
    .X(_0413_));
 sg13g2_nand2_2 _2922_ (.Y(_0783_),
    .A(_0722_),
    .B(_0781_));
 sg13g2_mux2_1 _2923_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .S(_0783_),
    .X(_0412_));
 sg13g2_mux2_1 _2924_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .S(_0783_),
    .X(_0411_));
 sg13g2_mux2_1 _2925_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ),
    .S(_0783_),
    .X(_0410_));
 sg13g2_mux2_1 _2926_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .S(_0783_),
    .X(_0409_));
 sg13g2_nand2_2 _2927_ (.Y(_0784_),
    .A(_0711_),
    .B(_0781_));
 sg13g2_mux2_1 _2928_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .S(_0784_),
    .X(_0408_));
 sg13g2_mux2_1 _2929_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .S(_0784_),
    .X(_0407_));
 sg13g2_mux2_1 _2930_ (.A0(net776),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .S(_0784_),
    .X(_0406_));
 sg13g2_mux2_1 _2931_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .S(_0784_),
    .X(_0405_));
 sg13g2_nor2_2 _2932_ (.A(_0714_),
    .B(_0728_),
    .Y(_0785_));
 sg13g2_mux2_1 _2933_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .A1(net753),
    .S(_0785_),
    .X(_0404_));
 sg13g2_mux2_1 _2934_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .A1(net762),
    .S(_0785_),
    .X(_0403_));
 sg13g2_mux2_1 _2935_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .A1(net773),
    .S(_0785_),
    .X(_0402_));
 sg13g2_mux2_1 _2936_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .A1(net784),
    .S(_0785_),
    .X(_0401_));
 sg13g2_nand2b_2 _2937_ (.Y(_0786_),
    .B(_0781_),
    .A_N(_0726_));
 sg13g2_mux2_1 _2938_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .S(_0786_),
    .X(_0400_));
 sg13g2_nor2_1 _2939_ (.A(net764),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_a21oi_1 _2940_ (.A1(_0634_),
    .A2(_0786_),
    .Y(_0399_),
    .B1(_0787_));
 sg13g2_nor2_1 _2941_ (.A(net776),
    .B(_0786_),
    .Y(_0788_));
 sg13g2_a21oi_1 _2942_ (.A1(_0635_),
    .A2(_0786_),
    .Y(_0398_),
    .B1(_0788_));
 sg13g2_nor2_1 _2943_ (.A(net787),
    .B(_0786_),
    .Y(_0789_));
 sg13g2_a21oi_1 _2944_ (.A1(_0636_),
    .A2(_0786_),
    .Y(_0397_),
    .B1(_0789_));
 sg13g2_nand2b_2 _2945_ (.Y(_0790_),
    .B(_0781_),
    .A_N(_0728_));
 sg13g2_mux2_1 _2946_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .S(_0790_),
    .X(_0396_));
 sg13g2_mux2_1 _2947_ (.A0(net765),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .S(_0790_),
    .X(_0395_));
 sg13g2_mux2_1 _2948_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .S(_0790_),
    .X(_0394_));
 sg13g2_mux2_1 _2949_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .S(_0790_),
    .X(_0393_));
 sg13g2_nand2b_2 _2950_ (.Y(_0791_),
    .B(_0781_),
    .A_N(_0707_));
 sg13g2_mux2_1 _2951_ (.A0(net755),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .S(_0791_),
    .X(_0392_));
 sg13g2_mux2_1 _2952_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .S(_0791_),
    .X(_0391_));
 sg13g2_mux2_1 _2953_ (.A0(net776),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .S(_0791_),
    .X(_0390_));
 sg13g2_mux2_1 _2954_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .S(_0791_),
    .X(_0389_));
 sg13g2_nor2_2 _2955_ (.A(_0719_),
    .B(_0737_),
    .Y(_0792_));
 sg13g2_mux2_1 _2956_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .A1(net760),
    .S(_0792_),
    .X(_0345_));
 sg13g2_mux2_1 _2957_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .A1(net770),
    .S(_0792_),
    .X(_0344_));
 sg13g2_mux2_1 _2958_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .A1(net782),
    .S(_0792_),
    .X(_0343_));
 sg13g2_mux2_1 _2959_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .A1(net793),
    .S(_0792_),
    .X(_0342_));
 sg13g2_nor2_2 _2960_ (.A(_0700_),
    .B(_0726_),
    .Y(_0793_));
 sg13g2_mux2_1 _2961_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .A1(net752),
    .S(_0793_),
    .X(_0341_));
 sg13g2_mux2_1 _2962_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .A1(net763),
    .S(_0793_),
    .X(_0340_));
 sg13g2_mux2_1 _2963_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .A1(net774),
    .S(_0793_),
    .X(_0339_));
 sg13g2_mux2_1 _2964_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .A1(net785),
    .S(_0793_),
    .X(_0338_));
 sg13g2_nand2b_2 _2965_ (.Y(_0794_),
    .B(_0732_),
    .A_N(_0728_));
 sg13g2_mux2_1 _2966_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .S(_0794_),
    .X(_0316_));
 sg13g2_mux2_1 _2967_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .S(_0794_),
    .X(_0315_));
 sg13g2_mux2_1 _2968_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .S(_0794_),
    .X(_0314_));
 sg13g2_mux2_1 _2969_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .S(_0794_),
    .X(_0313_));
 sg13g2_nand2b_2 _2970_ (.Y(_0795_),
    .B(_0720_),
    .A_N(_0714_));
 sg13g2_mux2_1 _2971_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .S(_0795_),
    .X(_0312_));
 sg13g2_mux2_1 _2972_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .S(_0795_),
    .X(_0311_));
 sg13g2_mux2_1 _2973_ (.A0(net775),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ),
    .S(_0795_),
    .X(_0310_));
 sg13g2_mux2_1 _2974_ (.A0(net786),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ),
    .S(_0795_),
    .X(_0309_));
 sg13g2_nand2_2 _2975_ (.Y(_0796_),
    .A(_0716_),
    .B(_0781_));
 sg13g2_nor2_1 _2976_ (.A(net754),
    .B(_0796_),
    .Y(_0797_));
 sg13g2_a21oi_1 _2977_ (.A1(_0649_),
    .A2(_0796_),
    .Y(_0298_),
    .B1(_0797_));
 sg13g2_mux2_1 _2978_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .S(_0796_),
    .X(_0297_));
 sg13g2_nor2_1 _2979_ (.A(net775),
    .B(_0796_),
    .Y(_0798_));
 sg13g2_a21oi_1 _2980_ (.A1(_0650_),
    .A2(_0796_),
    .Y(_0296_),
    .B1(_0798_));
 sg13g2_mux2_1 _2981_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .S(_0796_),
    .X(_0295_));
 sg13g2_nand2_2 _2982_ (.Y(_0799_),
    .A(_0699_),
    .B(_0722_));
 sg13g2_mux2_1 _2983_ (.A0(net753),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .S(_0799_),
    .X(_0294_));
 sg13g2_mux2_1 _2984_ (.A0(net762),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .S(_0799_),
    .X(_0293_));
 sg13g2_mux2_1 _2985_ (.A0(net773),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .S(_0799_),
    .X(_0292_));
 sg13g2_mux2_1 _2986_ (.A0(net784),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .S(_0799_),
    .X(_0291_));
 sg13g2_nand2_2 _2987_ (.Y(_0800_),
    .A(_0722_),
    .B(_0771_));
 sg13g2_mux2_1 _2988_ (.A0(net759),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .S(_0800_),
    .X(_0290_));
 sg13g2_mux2_1 _2989_ (.A0(net771),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .S(_0800_),
    .X(_0289_));
 sg13g2_mux2_1 _2990_ (.A0(net781),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .S(_0800_),
    .X(_0288_));
 sg13g2_mux2_1 _2991_ (.A0(net791),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ),
    .S(_0800_),
    .X(_0287_));
 sg13g2_nor2_2 _2992_ (.A(_0707_),
    .B(_0714_),
    .Y(_0801_));
 sg13g2_mux2_1 _2993_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .A1(net756),
    .S(_0801_),
    .X(_0286_));
 sg13g2_mux2_1 _2994_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .A1(net763),
    .S(_0801_),
    .X(_0285_));
 sg13g2_mux2_1 _2995_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .A1(net774),
    .S(_0801_),
    .X(_0284_));
 sg13g2_mux2_1 _2996_ (.A0(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .A1(net785),
    .S(_0801_),
    .X(_0283_));
 sg13g2_nand2b_2 _2997_ (.Y(_0802_),
    .B(_0781_),
    .A_N(_0737_));
 sg13g2_mux2_1 _2998_ (.A0(net754),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .S(_0802_),
    .X(_0282_));
 sg13g2_mux2_1 _2999_ (.A0(net764),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .S(_0802_),
    .X(_0281_));
 sg13g2_mux2_1 _3000_ (.A0(net776),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .S(_0802_),
    .X(_0280_));
 sg13g2_mux2_1 _3001_ (.A0(net787),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .S(_0802_),
    .X(_0279_));
 sg13g2_nand2_2 _3002_ (.Y(_0803_),
    .A(_0716_),
    .B(_0744_));
 sg13g2_mux2_1 _3003_ (.A0(net758),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .S(_0803_),
    .X(_0270_));
 sg13g2_mux2_1 _3004_ (.A0(net768),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .S(_0803_),
    .X(_0269_));
 sg13g2_mux2_1 _3005_ (.A0(net779),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .S(_0803_),
    .X(_0268_));
 sg13g2_mux2_1 _3006_ (.A0(net789),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .S(_0803_),
    .X(_0267_));
 sg13g2_and2_1 _3007_ (.A(net629),
    .B(_0680_),
    .X(_0804_));
 sg13g2_nand2_1 _3008_ (.Y(_0805_),
    .A(net629),
    .B(_0680_));
 sg13g2_and2_1 _3009_ (.A(\videogen.fancy_shader.video_x[8] ),
    .B(\videogen.fancy_shader.video_x[9] ),
    .X(_0806_));
 sg13g2_nor4_2 _3010_ (.A(\videogen.fancy_shader.video_y[9] ),
    .B(_0674_),
    .C(_0804_),
    .Y(_0807_),
    .D(_0806_));
 sg13g2_and2_1 _3011_ (.A(net795),
    .B(_0807_),
    .X(_0371_));
 sg13g2_nor2_2 _3012_ (.A(net746),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ),
    .Y(_0808_));
 sg13g2_nand2b_2 _3013_ (.Y(_0809_),
    .B(net795),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ));
 sg13g2_and2_1 _3014_ (.A(\videogen.fancy_shader.video_x[1] ),
    .B(\videogen.fancy_shader.video_x[0] ),
    .X(_0810_));
 sg13g2_and2_1 _3015_ (.A(\videogen.fancy_shader.video_x[2] ),
    .B(_0810_),
    .X(_0811_));
 sg13g2_and2_1 _3016_ (.A(\videogen.fancy_shader.video_x[3] ),
    .B(_0811_),
    .X(_0812_));
 sg13g2_nand2_1 _3017_ (.Y(_0813_),
    .A(\videogen.fancy_shader.video_x[3] ),
    .B(_0811_));
 sg13g2_and2_1 _3018_ (.A(\videogen.fancy_shader.video_x[4] ),
    .B(_0812_),
    .X(_0814_));
 sg13g2_and2_1 _3019_ (.A(\videogen.fancy_shader.video_x[5] ),
    .B(_0814_),
    .X(_0815_));
 sg13g2_and2_1 _3020_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(_0815_),
    .X(_0816_));
 sg13g2_and2_1 _3021_ (.A(_0651_),
    .B(_0680_),
    .X(_0817_));
 sg13g2_and2_1 _3022_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .B(_0807_),
    .X(_0818_));
 sg13g2_nand3_1 _3023_ (.B(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .Y(_0819_));
 sg13g2_or2_1 _3024_ (.X(_0820_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ));
 sg13g2_nor4_1 _3025_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .C(_0819_),
    .D(_0820_),
    .Y(_0821_));
 sg13g2_a22oi_1 _3026_ (.Y(_0822_),
    .B1(_0818_),
    .B2(_0821_),
    .A2(_0817_),
    .A1(_0816_));
 sg13g2_nand2b_1 _3027_ (.Y(_0823_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ),
    .A_N(_0807_));
 sg13g2_or2_1 _3028_ (.X(_0824_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.state[3] ),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ));
 sg13g2_nand2_1 _3029_ (.Y(_0825_),
    .A(net796),
    .B(_0824_));
 sg13g2_nand4_1 _3030_ (.B(_0822_),
    .C(_0823_),
    .A(net795),
    .Y(_0826_),
    .D(_0824_));
 sg13g2_a21oi_1 _3031_ (.A1(_0808_),
    .A2(_0826_),
    .Y(_0002_),
    .B1(_0371_));
 sg13g2_o21ai_1 _3032_ (.B1(_0807_),
    .Y(_0827_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ),
    .A2(_0822_));
 sg13g2_a21oi_1 _3033_ (.A1(_0659_),
    .A2(_0827_),
    .Y(_0003_),
    .B1(net746));
 sg13g2_nor3_1 _3034_ (.A(\serialize.bit_cnt[1] ),
    .B(net412),
    .C(net415),
    .Y(\serialize.n410 ));
 sg13g2_a21oi_2 _3035_ (.B1(net595),
    .Y(net8),
    .A2(net549),
    .A1(net628));
 sg13g2_a21oi_1 _3036_ (.A1(net549),
    .A2(_0703_),
    .Y(net9),
    .B1(net595));
 sg13g2_a21oi_2 _3037_ (.B1(net595),
    .Y(net10),
    .A2(_0709_),
    .A1(net549));
 sg13g2_a21oi_2 _3038_ (.B1(net595),
    .Y(net11),
    .A2(_0690_),
    .A1(net549));
 sg13g2_a21oi_2 _3039_ (.B1(net595),
    .Y(net12),
    .A2(_0693_),
    .A1(net549));
 sg13g2_a21oi_2 _3040_ (.B1(net595),
    .Y(net13),
    .A2(_0695_),
    .A1(net549));
 sg13g2_nor2_1 _3041_ (.A(_0683_),
    .B(_0694_),
    .Y(_0828_));
 sg13g2_nand2_1 _3042_ (.Y(_0829_),
    .A(\videogen.fancy_shader.video_y[3] ),
    .B(\videogen.fancy_shader.video_y[2] ));
 sg13g2_nand2b_1 _3043_ (.Y(_0830_),
    .B(\videogen.fancy_shader.video_y[4] ),
    .A_N(\videogen.fancy_shader.video_y[5] ));
 sg13g2_nand2_1 _3044_ (.Y(_0831_),
    .A(\videogen.fancy_shader.video_y[1] ),
    .B(net608));
 sg13g2_nand4_1 _3045_ (.B(\videogen.fancy_shader.video_y[8] ),
    .C(\videogen.fancy_shader.video_y[7] ),
    .A(_0637_),
    .Y(_0832_),
    .D(\videogen.fancy_shader.video_y[6] ));
 sg13g2_nor4_1 _3046_ (.A(_0829_),
    .B(_0830_),
    .C(_0831_),
    .D(_0832_),
    .Y(_0833_));
 sg13g2_nor2_1 _3047_ (.A(_0829_),
    .B(_0831_),
    .Y(_0834_));
 sg13g2_nor2_2 _3048_ (.A(_0677_),
    .B(_0833_),
    .Y(_0835_));
 sg13g2_o21ai_1 _3049_ (.B1(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .Y(_0836_),
    .A1(_0828_),
    .A2(_0835_));
 sg13g2_nand3_1 _3050_ (.B(net549),
    .C(_0694_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .Y(_0837_));
 sg13g2_a21o_1 _3051_ (.A2(_0694_),
    .A1(net549),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .X(_0838_));
 sg13g2_nand2_1 _3052_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_a21oi_1 _3053_ (.A1(_0835_),
    .A2(_0839_),
    .Y(net14),
    .B1(_0836_));
 sg13g2_nor2_2 _3054_ (.A(_0648_),
    .B(_0837_),
    .Y(_0840_));
 sg13g2_xnor2_1 _3055_ (.Y(_0841_),
    .A(_0648_),
    .B(_0837_));
 sg13g2_a21oi_1 _3056_ (.A1(_0835_),
    .A2(_0841_),
    .Y(net15),
    .B1(_0836_));
 sg13g2_xnor2_1 _3057_ (.Y(_0842_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(_0840_));
 sg13g2_a21oi_1 _3058_ (.A1(_0835_),
    .A2(_0842_),
    .Y(net16),
    .B1(_0836_));
 sg13g2_nand3_1 _3059_ (.B(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .C(_0840_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .Y(_0843_));
 sg13g2_a21o_1 _3060_ (.A2(_0840_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .X(_0844_));
 sg13g2_nand2_1 _3061_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_a21oi_1 _3062_ (.A1(_0835_),
    .A2(_0845_),
    .Y(net17),
    .B1(_0836_));
 sg13g2_nand4_1 _3063_ (.B(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .Y(_0846_),
    .D(_0840_));
 sg13g2_xor2_1 _3064_ (.B(_0843_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .X(_0847_));
 sg13g2_a21oi_1 _3065_ (.A1(_0835_),
    .A2(_0847_),
    .Y(net18),
    .B1(_0836_));
 sg13g2_o21ai_1 _3066_ (.B1(_0835_),
    .Y(_0848_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0846_));
 sg13g2_a21oi_1 _3067_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0846_),
    .Y(_0849_),
    .B1(_0848_));
 sg13g2_nor2_1 _3068_ (.A(_0836_),
    .B(_0849_),
    .Y(net7));
 sg13g2_mux2_1 _3069_ (.A0(\serialize.n461 ),
    .A1(\serialize.n459 ),
    .S(clknet_1_0__leaf_clk),
    .X(net4));
 sg13g2_mux2_1 _3070_ (.A0(\serialize.n458 ),
    .A1(\serialize.n456 ),
    .S(clknet_1_0__leaf_clk),
    .X(net3));
 sg13g2_mux2_1 _3071_ (.A0(\serialize.n455 ),
    .A1(\serialize.n453 ),
    .S(clknet_1_1__leaf_clk),
    .X(net5));
 sg13g2_mux2_1 _3072_ (.A0(\serialize.n452 ),
    .A1(\serialize.n450 ),
    .S(clknet_1_1__leaf_clk),
    .X(net6));
 sg13g2_nor2_1 _3073_ (.A(net412),
    .B(net695),
    .Y(\serialize.n433[0] ));
 sg13g2_nor2b_1 _3074_ (.A(net697),
    .B_N(net410),
    .Y(\serialize.n431[0] ));
 sg13g2_nor2b_1 _3075_ (.A(net697),
    .B_N(net411),
    .Y(\serialize.n431[1] ));
 sg13g2_nor2b_1 _3076_ (.A(net697),
    .B_N(net408),
    .Y(\serialize.n431[2] ));
 sg13g2_nor2b_1 _3077_ (.A(net697),
    .B_N(net409),
    .Y(\serialize.n431[3] ));
 sg13g2_nor2b_1 _3078_ (.A(net697),
    .B_N(net413),
    .Y(\serialize.n431[4] ));
 sg13g2_or2_1 _3079_ (.X(\serialize.n431[5] ),
    .B(net697),
    .A(net413));
 sg13g2_or2_1 _3080_ (.X(\serialize.n431[6] ),
    .B(net700),
    .A(net419));
 sg13g2_mux2_1 _3081_ (.A0(net428),
    .A1(\blue_tmds_par[0] ),
    .S(net697),
    .X(\serialize.n429[0] ));
 sg13g2_mux2_1 _3082_ (.A0(net440),
    .A1(\blue_tmds_par[1] ),
    .S(net694),
    .X(\serialize.n429[1] ));
 sg13g2_mux2_1 _3083_ (.A0(net437),
    .A1(\blue_tmds_par[2] ),
    .S(net694),
    .X(\serialize.n429[2] ));
 sg13g2_mux2_1 _3084_ (.A0(net433),
    .A1(\blue_tmds_par[3] ),
    .S(net700),
    .X(\serialize.n429[3] ));
 sg13g2_mux2_1 _3085_ (.A0(net443),
    .A1(\blue_tmds_par[2] ),
    .S(net700),
    .X(\serialize.n429[4] ));
 sg13g2_mux2_1 _3086_ (.A0(net427),
    .A1(\blue_tmds_par[5] ),
    .S(net694),
    .X(\serialize.n429[5] ));
 sg13g2_mux2_1 _3087_ (.A0(net435),
    .A1(\blue_tmds_par[6] ),
    .S(net694),
    .X(\serialize.n429[6] ));
 sg13g2_mux2_1 _3088_ (.A0(net425),
    .A1(\blue_tmds_par[7] ),
    .S(net694),
    .X(\serialize.n429[7] ));
 sg13g2_and2_1 _3089_ (.A(\blue_tmds_par[8] ),
    .B(net694),
    .X(\serialize.n429[8] ));
 sg13g2_and2_1 _3090_ (.A(\blue_tmds_par[9] ),
    .B(net694),
    .X(\serialize.n429[9] ));
 sg13g2_mux2_1 _3091_ (.A0(net423),
    .A1(\green_tmds_par[0] ),
    .S(net696),
    .X(\serialize.n428[0] ));
 sg13g2_nand2_1 _3092_ (.Y(_0850_),
    .A(\green_tmds_par[1] ),
    .B(net698));
 sg13g2_o21ai_1 _3093_ (.B1(_0850_),
    .Y(\serialize.n428[1] ),
    .A1(_0668_),
    .A2(net696));
 sg13g2_mux2_1 _3094_ (.A0(net436),
    .A1(\green_tmds_par[2] ),
    .S(net696),
    .X(\serialize.n428[2] ));
 sg13g2_o21ai_1 _3095_ (.B1(_0850_),
    .Y(\serialize.n428[3] ),
    .A1(_0669_),
    .A2(net698));
 sg13g2_mux2_1 _3096_ (.A0(net439),
    .A1(\green_tmds_par[2] ),
    .S(net695),
    .X(\serialize.n428[4] ));
 sg13g2_o21ai_1 _3097_ (.B1(_0850_),
    .Y(\serialize.n428[5] ),
    .A1(_0670_),
    .A2(net698));
 sg13g2_mux2_1 _3098_ (.A0(net429),
    .A1(\green_tmds_par[6] ),
    .S(net695),
    .X(\serialize.n428[6] ));
 sg13g2_mux2_1 _3099_ (.A0(net438),
    .A1(\green_tmds_par[7] ),
    .S(net698),
    .X(\serialize.n428[7] ));
 sg13g2_and2_1 _3100_ (.A(\green_tmds_par[8] ),
    .B(net695),
    .X(\serialize.n428[8] ));
 sg13g2_and2_1 _3101_ (.A(\green_tmds_par[9] ),
    .B(net697),
    .X(\serialize.n428[9] ));
 sg13g2_mux2_1 _3102_ (.A0(net421),
    .A1(\red_tmds_par[0] ),
    .S(net699),
    .X(\serialize.n427[0] ));
 sg13g2_mux2_1 _3103_ (.A0(net441),
    .A1(\red_tmds_par[1] ),
    .S(net699),
    .X(\serialize.n427[1] ));
 sg13g2_mux2_1 _3104_ (.A0(net422),
    .A1(\red_tmds_par[2] ),
    .S(net696),
    .X(\serialize.n427[2] ));
 sg13g2_mux2_1 _3105_ (.A0(net424),
    .A1(\red_tmds_par[3] ),
    .S(net696),
    .X(\serialize.n427[3] ));
 sg13g2_mux2_1 _3106_ (.A0(net442),
    .A1(\red_tmds_par[4] ),
    .S(net696),
    .X(\serialize.n427[4] ));
 sg13g2_mux2_1 _3107_ (.A0(net426),
    .A1(\red_tmds_par[5] ),
    .S(net696),
    .X(\serialize.n427[5] ));
 sg13g2_mux2_1 _3108_ (.A0(net430),
    .A1(\red_tmds_par[6] ),
    .S(net695),
    .X(\serialize.n427[6] ));
 sg13g2_mux2_1 _3109_ (.A0(net431),
    .A1(\red_tmds_par[7] ),
    .S(net696),
    .X(\serialize.n427[7] ));
 sg13g2_and2_1 _3110_ (.A(\red_tmds_par[8] ),
    .B(net695),
    .X(\serialize.n427[8] ));
 sg13g2_and2_1 _3111_ (.A(\red_tmds_par[9] ),
    .B(net695),
    .X(\serialize.n427[9] ));
 sg13g2_nor2_1 _3112_ (.A(net677),
    .B(net729),
    .Y(_0006_));
 sg13g2_inv_1 _3113_ (.Y(clk_video),
    .A(_0006_));
 sg13g2_nand2_1 _3114_ (.Y(_0851_),
    .A(net795),
    .B(_0822_));
 sg13g2_nor2_1 _3115_ (.A(_0823_),
    .B(_0851_),
    .Y(_0001_));
 sg13g2_nor2_1 _3116_ (.A(_0822_),
    .B(_0825_),
    .Y(_0000_));
 sg13g2_and2_1 _3117_ (.A(net606),
    .B(net803),
    .X(_0852_));
 sg13g2_nand2_1 _3118_ (.Y(_0853_),
    .A(net607),
    .B(net799));
 sg13g2_and2_1 _3119_ (.A(\tmds_green.dc_balancing_reg[0] ),
    .B(_0852_),
    .X(_0263_));
 sg13g2_and2_1 _3120_ (.A(\tmds_blue.dc_balancing_reg[0] ),
    .B(_0852_),
    .X(_0264_));
 sg13g2_o21ai_1 _3121_ (.B1(net796),
    .Y(_0854_),
    .A1(net739),
    .A2(net432));
 sg13g2_a21oi_1 _3122_ (.A1(net739),
    .A2(net432),
    .Y(_0265_),
    .B1(_0854_));
 sg13g2_and3_1 _3123_ (.X(_0266_),
    .A(net796),
    .B(net739),
    .C(net432));
 sg13g2_nor2_1 _3124_ (.A(_0654_),
    .B(net571),
    .Y(_0271_));
 sg13g2_nor4_1 _3125_ (.A(\tmds_green.dc_balancing_reg[0] ),
    .B(\tmds_green.dc_balancing_reg[1] ),
    .C(\tmds_green.dc_balancing_reg[3] ),
    .D(\tmds_green.dc_balancing_reg[2] ),
    .Y(_0855_));
 sg13g2_and2_1 _3126_ (.A(_0654_),
    .B(_0855_),
    .X(_0856_));
 sg13g2_nand2b_1 _3127_ (.Y(_0857_),
    .B(net600),
    .A_N(\tmds_green.n132 ));
 sg13g2_xor2_1 _3128_ (.B(net599),
    .A(net601),
    .X(_0858_));
 sg13g2_nand2_1 _3129_ (.Y(_0859_),
    .A(\tmds_green.n100 ),
    .B(_0654_));
 sg13g2_nand2_1 _3130_ (.Y(_0860_),
    .A(net601),
    .B(_0856_));
 sg13g2_mux2_1 _3131_ (.A0(_0858_),
    .A1(net599),
    .S(_0856_),
    .X(_0861_));
 sg13g2_nand2b_1 _3132_ (.Y(_0862_),
    .B(\tmds_green.dc_balancing_reg[4] ),
    .A_N(net601));
 sg13g2_o21ai_1 _3133_ (.B1(_0862_),
    .Y(_0863_),
    .A1(_0855_),
    .A2(_0859_));
 sg13g2_xor2_1 _3134_ (.B(_0863_),
    .A(\tmds_green.n126 ),
    .X(_0864_));
 sg13g2_o21ai_1 _3135_ (.B1(_0852_),
    .Y(_0865_),
    .A1(_0861_),
    .A2(_0864_));
 sg13g2_a21oi_1 _3136_ (.A1(_0861_),
    .A2(_0864_),
    .Y(_0273_),
    .B1(_0865_));
 sg13g2_nor4_1 _3137_ (.A(\tmds_red.dc_balancing_reg[1] ),
    .B(\tmds_red.dc_balancing_reg[0] ),
    .C(\tmds_red.dc_balancing_reg[3] ),
    .D(\tmds_red.dc_balancing_reg[2] ),
    .Y(_0866_));
 sg13g2_nand2_1 _3138_ (.Y(_0867_),
    .A(\tmds_red.n114 ),
    .B(\tmds_red.n132 ));
 sg13g2_nor2_1 _3139_ (.A(\tmds_red.n114 ),
    .B(\tmds_red.n132 ),
    .Y(_0868_));
 sg13g2_xnor2_1 _3140_ (.Y(_0869_),
    .A(\tmds_red.n114 ),
    .B(\tmds_red.n132 ));
 sg13g2_a21oi_1 _3141_ (.A1(\tmds_red.n126 ),
    .A2(\tmds_red.n132 ),
    .Y(_0870_),
    .B1(\tmds_red.n100 ));
 sg13g2_nor2_1 _3142_ (.A(\tmds_red.n126 ),
    .B(\tmds_red.n132 ),
    .Y(_0871_));
 sg13g2_nor2_1 _3143_ (.A(_0870_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_xnor2_1 _3144_ (.Y(_0873_),
    .A(\tmds_red.n114 ),
    .B(_0872_));
 sg13g2_xor2_1 _3145_ (.B(\tmds_red.n132 ),
    .A(\tmds_red.n126 ),
    .X(_0874_));
 sg13g2_xnor2_1 _3146_ (.Y(_0875_),
    .A(\tmds_red.n100 ),
    .B(_0874_));
 sg13g2_nor3_1 _3147_ (.A(_0663_),
    .B(_0873_),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_nand2b_1 _3148_ (.Y(_0877_),
    .B(\tmds_red.n114 ),
    .A_N(_0870_));
 sg13g2_xnor2_1 _3149_ (.Y(_0878_),
    .A(_0876_),
    .B(_0877_));
 sg13g2_nand2_1 _3150_ (.Y(_0879_),
    .A(_0663_),
    .B(_0875_));
 sg13g2_xor2_1 _3151_ (.B(_0879_),
    .A(_0873_),
    .X(_0880_));
 sg13g2_a21oi_1 _3152_ (.A1(\tmds_red.n100 ),
    .A2(_0880_),
    .Y(_0881_),
    .B1(_0878_));
 sg13g2_xnor2_1 _3153_ (.Y(_0882_),
    .A(\tmds_red.n100 ),
    .B(\tmds_red.n102 ));
 sg13g2_xor2_1 _3154_ (.B(_0882_),
    .A(net547),
    .X(_0883_));
 sg13g2_inv_1 _3155_ (.Y(_0884_),
    .A(_0883_));
 sg13g2_xnor2_1 _3156_ (.Y(_0885_),
    .A(_0869_),
    .B(_0883_));
 sg13g2_nor2_1 _3157_ (.A(\tmds_red.n102 ),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_nor2_1 _3158_ (.A(net548),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_nand2_1 _3159_ (.Y(_0888_),
    .A(\tmds_red.n100 ),
    .B(_0869_));
 sg13g2_a21oi_1 _3160_ (.A1(_0867_),
    .A2(_0882_),
    .Y(_0889_),
    .B1(_0868_));
 sg13g2_nand2b_1 _3161_ (.Y(_0890_),
    .B(\tmds_red.n126 ),
    .A_N(\tmds_red.n132 ));
 sg13g2_o21ai_1 _3162_ (.B1(_0890_),
    .Y(_0891_),
    .A1(_0874_),
    .A2(net547));
 sg13g2_xnor2_1 _3163_ (.Y(_0892_),
    .A(_0889_),
    .B(_0891_));
 sg13g2_inv_1 _3164_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_xnor2_1 _3165_ (.Y(_0894_),
    .A(_0869_),
    .B(_0892_));
 sg13g2_nand2_1 _3166_ (.Y(_0895_),
    .A(_0883_),
    .B(_0894_));
 sg13g2_o21ai_1 _3167_ (.B1(_0895_),
    .Y(_0896_),
    .A1(_0883_),
    .A2(_0893_));
 sg13g2_a21oi_1 _3168_ (.A1(\tmds_red.n102 ),
    .A2(_0885_),
    .Y(_0897_),
    .B1(_0887_));
 sg13g2_xor2_1 _3169_ (.B(_0897_),
    .A(_0896_),
    .X(_0898_));
 sg13g2_nand2b_1 _3170_ (.Y(_0899_),
    .B(_0898_),
    .A_N(_0888_));
 sg13g2_a22oi_1 _3171_ (.Y(_0900_),
    .B1(_0895_),
    .B2(_0897_),
    .A2(_0892_),
    .A1(_0884_));
 sg13g2_nor2b_2 _3172_ (.A(_0900_),
    .B_N(_0899_),
    .Y(_0901_));
 sg13g2_nor2b_2 _3173_ (.A(_0899_),
    .B_N(_0900_),
    .Y(_0902_));
 sg13g2_nor2_1 _3174_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_xor2_1 _3175_ (.B(_0898_),
    .A(_0888_),
    .X(_0904_));
 sg13g2_and2_1 _3176_ (.A(_0869_),
    .B(_0904_),
    .X(_0905_));
 sg13g2_a22oi_1 _3177_ (.Y(_0906_),
    .B1(_0903_),
    .B2(_0905_),
    .A2(_0866_),
    .A1(_0664_));
 sg13g2_nand2b_1 _3178_ (.Y(_0907_),
    .B(_0903_),
    .A_N(_0905_));
 sg13g2_nand2b_1 _3179_ (.Y(_0908_),
    .B(_0907_),
    .A_N(_0902_));
 sg13g2_nor2_1 _3180_ (.A(\tmds_red.dc_balancing_reg[4] ),
    .B(_0866_),
    .Y(_0909_));
 sg13g2_a22oi_1 _3181_ (.Y(_0910_),
    .B1(_0908_),
    .B2(_0909_),
    .A2(_0901_),
    .A1(\tmds_red.dc_balancing_reg[4] ));
 sg13g2_nand2_1 _3182_ (.Y(_0911_),
    .A(_0906_),
    .B(_0910_));
 sg13g2_inv_1 _3183_ (.Y(_0912_),
    .A(_0911_));
 sg13g2_nor2b_2 _3184_ (.A(_0906_),
    .B_N(net547),
    .Y(_0913_));
 sg13g2_nor2_2 _3185_ (.A(_0912_),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_o21ai_1 _3186_ (.B1(_0852_),
    .Y(_0915_),
    .A1(\tmds_red.n100 ),
    .A2(_0914_));
 sg13g2_a21oi_1 _3187_ (.A1(\tmds_red.n100 ),
    .A2(_0914_),
    .Y(_0274_),
    .B1(_0915_));
 sg13g2_nand2_1 _3188_ (.Y(_0916_),
    .A(net547),
    .B(_0910_));
 sg13g2_o21ai_1 _3189_ (.B1(_0916_),
    .Y(_0917_),
    .A1(net547),
    .A2(_0912_));
 sg13g2_nor2_1 _3190_ (.A(net571),
    .B(_0917_),
    .Y(_0275_));
 sg13g2_o21ai_1 _3191_ (.B1(_0852_),
    .Y(_0918_),
    .A1(_0882_),
    .A2(_0917_));
 sg13g2_a21oi_1 _3192_ (.A1(_0882_),
    .A2(_0917_),
    .Y(_0276_),
    .B1(_0918_));
 sg13g2_xnor2_1 _3193_ (.Y(_0919_),
    .A(_0663_),
    .B(_0875_));
 sg13g2_o21ai_1 _3194_ (.B1(_0852_),
    .Y(_0920_),
    .A1(_0917_),
    .A2(_0919_));
 sg13g2_a21oi_1 _3195_ (.A1(_0917_),
    .A2(_0919_),
    .Y(_0278_),
    .B1(_0920_));
 sg13g2_nor3_1 _3196_ (.A(net629),
    .B(\videogen.fancy_shader.video_x[6] ),
    .C(\videogen.fancy_shader.video_x[5] ),
    .Y(_0921_));
 sg13g2_and3_2 _3197_ (.X(_0922_),
    .A(_0806_),
    .B(_0814_),
    .C(_0921_));
 sg13g2_nand2b_2 _3198_ (.Y(_0923_),
    .B(net797),
    .A_N(_0922_));
 sg13g2_nor2_1 _3199_ (.A(\videogen.fancy_shader.video_x[0] ),
    .B(_0923_),
    .Y(_0299_));
 sg13g2_nor3_1 _3200_ (.A(_0681_),
    .B(_0810_),
    .C(_0923_),
    .Y(_0300_));
 sg13g2_nor2_1 _3201_ (.A(\videogen.fancy_shader.video_x[2] ),
    .B(_0810_),
    .Y(_0924_));
 sg13g2_nor3_1 _3202_ (.A(net750),
    .B(_0811_),
    .C(_0924_),
    .Y(_0301_));
 sg13g2_o21ai_1 _3203_ (.B1(net797),
    .Y(_0925_),
    .A1(\videogen.fancy_shader.video_x[3] ),
    .A2(_0811_));
 sg13g2_nor2_1 _3204_ (.A(_0812_),
    .B(_0925_),
    .Y(_0302_));
 sg13g2_nand2b_1 _3205_ (.Y(_0926_),
    .B(_0813_),
    .A_N(\videogen.fancy_shader.video_x[4] ));
 sg13g2_nand2_1 _3206_ (.Y(_0927_),
    .A(net797),
    .B(_0926_));
 sg13g2_nor2_1 _3207_ (.A(_0814_),
    .B(_0927_),
    .Y(_0303_));
 sg13g2_nor2_1 _3208_ (.A(\videogen.fancy_shader.video_x[5] ),
    .B(_0814_),
    .Y(_0928_));
 sg13g2_nor3_1 _3209_ (.A(_0815_),
    .B(_0923_),
    .C(_0928_),
    .Y(_0304_));
 sg13g2_nor2_1 _3210_ (.A(\videogen.fancy_shader.video_x[6] ),
    .B(_0815_),
    .Y(_0929_));
 sg13g2_nor3_1 _3211_ (.A(_0816_),
    .B(_0923_),
    .C(_0929_),
    .Y(_0305_));
 sg13g2_and2_1 _3212_ (.A(net629),
    .B(_0816_),
    .X(_0930_));
 sg13g2_nor2_1 _3213_ (.A(net629),
    .B(_0816_),
    .Y(_0931_));
 sg13g2_nor3_1 _3214_ (.A(_0923_),
    .B(_0930_),
    .C(_0931_),
    .Y(_0306_));
 sg13g2_nand2_1 _3215_ (.Y(_0932_),
    .A(\videogen.fancy_shader.video_x[8] ),
    .B(_0930_));
 sg13g2_xnor2_1 _3216_ (.Y(_0933_),
    .A(\videogen.fancy_shader.video_x[8] ),
    .B(_0930_));
 sg13g2_nor2_1 _3217_ (.A(_0923_),
    .B(_0933_),
    .Y(_0307_));
 sg13g2_xor2_1 _3218_ (.B(_0932_),
    .A(\videogen.fancy_shader.video_x[9] ),
    .X(_0934_));
 sg13g2_nor2_1 _3219_ (.A(_0923_),
    .B(_0934_),
    .Y(_0308_));
 sg13g2_nand2_1 _3220_ (.Y(_0935_),
    .A(\videogen.fancy_shader.video_y[3] ),
    .B(_0640_));
 sg13g2_xnor2_1 _3221_ (.Y(_0936_),
    .A(\videogen.fancy_shader.video_y[1] ),
    .B(net608));
 sg13g2_nor2_1 _3222_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_a21oi_1 _3223_ (.A1(_0675_),
    .A2(_0937_),
    .Y(_0317_),
    .B1(net745));
 sg13g2_o21ai_1 _3224_ (.B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .Y(_0938_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .A2(_0820_));
 sg13g2_o21ai_1 _3225_ (.B1(_0684_),
    .Y(_0939_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .A2(_0824_));
 sg13g2_nor2_2 _3226_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_and2_1 _3227_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0940_),
    .X(_0941_));
 sg13g2_nand2_2 _3228_ (.Y(_0942_),
    .A(_0677_),
    .B(_0683_));
 sg13g2_nand2_2 _3229_ (.Y(_0943_),
    .A(net796),
    .B(_0942_));
 sg13g2_nor2_1 _3230_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .B(_0940_),
    .Y(_0944_));
 sg13g2_nor3_1 _3231_ (.A(_0941_),
    .B(_0943_),
    .C(_0944_),
    .Y(_0318_));
 sg13g2_nor2_1 _3232_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .B(_0941_),
    .Y(_0945_));
 sg13g2_and2_1 _3233_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .B(_0941_),
    .X(_0946_));
 sg13g2_nor3_1 _3234_ (.A(_0943_),
    .B(_0945_),
    .C(_0946_),
    .Y(_0319_));
 sg13g2_nor2_1 _3235_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_and2_1 _3236_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .B(_0946_),
    .X(_0948_));
 sg13g2_nor3_1 _3237_ (.A(_0943_),
    .B(_0947_),
    .C(_0948_),
    .Y(_0320_));
 sg13g2_nor2_1 _3238_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_and2_1 _3239_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .B(_0948_),
    .X(_0950_));
 sg13g2_nor3_1 _3240_ (.A(_0943_),
    .B(_0949_),
    .C(_0950_),
    .Y(_0321_));
 sg13g2_nor2_1 _3241_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_and2_1 _3242_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .B(_0950_),
    .X(_0952_));
 sg13g2_nor3_1 _3243_ (.A(_0943_),
    .B(_0951_),
    .C(_0952_),
    .Y(_0322_));
 sg13g2_a21oi_1 _3244_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0952_),
    .Y(_0953_),
    .B1(_0943_));
 sg13g2_o21ai_1 _3245_ (.B1(_0953_),
    .Y(_0954_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .A2(_0952_));
 sg13g2_inv_1 _3246_ (.Y(_0323_),
    .A(_0954_));
 sg13g2_or3_1 _3247_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .C(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .X(_0955_));
 sg13g2_nand3_1 _3248_ (.B(_0807_),
    .C(_0955_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .Y(_0956_));
 sg13g2_inv_1 _3249_ (.Y(_0957_),
    .A(_0956_));
 sg13g2_o21ai_1 _3250_ (.B1(_0808_),
    .Y(_0958_),
    .A1(_0647_),
    .A2(_0956_));
 sg13g2_a21oi_1 _3251_ (.A1(_0647_),
    .A2(_0956_),
    .Y(_0324_),
    .B1(_0958_));
 sg13g2_nor2_1 _3252_ (.A(net578),
    .B(_0956_),
    .Y(_0959_));
 sg13g2_a21oi_1 _3253_ (.A1(net628),
    .A2(_0957_),
    .Y(_0960_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ));
 sg13g2_nor3_1 _3254_ (.A(_0809_),
    .B(_0959_),
    .C(_0960_),
    .Y(_0325_));
 sg13g2_xnor2_1 _3255_ (.Y(_0961_),
    .A(net623),
    .B(_0959_));
 sg13g2_nor2_1 _3256_ (.A(_0809_),
    .B(_0961_),
    .Y(_0326_));
 sg13g2_a21oi_1 _3257_ (.A1(net623),
    .A2(_0959_),
    .Y(_0962_),
    .B1(net616));
 sg13g2_nor4_1 _3258_ (.A(net596),
    .B(_0646_),
    .C(net578),
    .D(_0956_),
    .Y(_0963_));
 sg13g2_nor3_1 _3259_ (.A(_0809_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0327_));
 sg13g2_or2_1 _3260_ (.X(_0964_),
    .B(_0963_),
    .A(net611));
 sg13g2_nand2_1 _3261_ (.Y(_0965_),
    .A(net611),
    .B(_0963_));
 sg13g2_and3_1 _3262_ (.X(_0328_),
    .A(_0808_),
    .B(_0964_),
    .C(_0965_));
 sg13g2_xor2_1 _3263_ (.B(_0965_),
    .A(net610),
    .X(_0966_));
 sg13g2_nor2_1 _3264_ (.A(_0809_),
    .B(_0966_),
    .Y(_0329_));
 sg13g2_or2_1 _3265_ (.X(_0967_),
    .B(_0943_),
    .A(_0940_));
 sg13g2_nor2b_1 _3266_ (.A(_0939_),
    .B_N(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .Y(_0968_));
 sg13g2_nor2b_1 _3267_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .B_N(_0939_),
    .Y(_0969_));
 sg13g2_nor3_1 _3268_ (.A(_0967_),
    .B(_0968_),
    .C(_0969_),
    .Y(_0330_));
 sg13g2_nor2_1 _3269_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .B(_0968_),
    .Y(_0970_));
 sg13g2_and2_1 _3270_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .B(_0968_),
    .X(_0971_));
 sg13g2_nor3_1 _3271_ (.A(_0967_),
    .B(_0970_),
    .C(_0971_),
    .Y(_0331_));
 sg13g2_a21oi_1 _3272_ (.A1(_0938_),
    .A2(_0971_),
    .Y(_0972_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ));
 sg13g2_and2_1 _3273_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .B(_0971_),
    .X(_0973_));
 sg13g2_nor3_1 _3274_ (.A(_0967_),
    .B(_0972_),
    .C(_0973_),
    .Y(_0332_));
 sg13g2_nor2_1 _3275_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_nor2_1 _3276_ (.A(_0967_),
    .B(_0974_),
    .Y(_0333_));
 sg13g2_nand2_2 _3277_ (.Y(_0975_),
    .A(_0808_),
    .B(_0956_));
 sg13g2_nor2_1 _3278_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .B(_0807_),
    .Y(_0976_));
 sg13g2_nor3_1 _3279_ (.A(_0818_),
    .B(_0975_),
    .C(_0976_),
    .Y(_0334_));
 sg13g2_and2_1 _3280_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .B(_0818_),
    .X(_0977_));
 sg13g2_nor2_1 _3281_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .B(_0818_),
    .Y(_0978_));
 sg13g2_nor3_1 _3282_ (.A(_0975_),
    .B(_0977_),
    .C(_0978_),
    .Y(_0335_));
 sg13g2_xnor2_1 _3283_ (.Y(_0979_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .B(_0977_));
 sg13g2_nor2_1 _3284_ (.A(_0975_),
    .B(_0979_),
    .Y(_0336_));
 sg13g2_a21oi_1 _3285_ (.A1(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .A2(_0977_),
    .Y(_0980_),
    .B1(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ));
 sg13g2_nor2_1 _3286_ (.A(_0975_),
    .B(_0980_),
    .Y(_0337_));
 sg13g2_nor2_2 _3287_ (.A(_0643_),
    .B(_0942_),
    .Y(_0981_));
 sg13g2_a21oi_1 _3288_ (.A1(_0643_),
    .A2(_0942_),
    .Y(_0982_),
    .B1(net750));
 sg13g2_nor2b_1 _3289_ (.A(_0981_),
    .B_N(_0982_),
    .Y(_0346_));
 sg13g2_o21ai_1 _3290_ (.B1(net798),
    .Y(_0983_),
    .A1(\videogen.fancy_shader.n646[1] ),
    .A2(_0981_));
 sg13g2_a21oi_1 _3291_ (.A1(\videogen.fancy_shader.n646[1] ),
    .A2(_0981_),
    .Y(_0347_),
    .B1(_0983_));
 sg13g2_a21oi_1 _3292_ (.A1(\videogen.fancy_shader.n646[1] ),
    .A2(_0981_),
    .Y(_0984_),
    .B1(\videogen.fancy_shader.n646[2] ));
 sg13g2_nand2_1 _3293_ (.Y(_0985_),
    .A(\videogen.fancy_shader.video_y[1] ),
    .B(\videogen.fancy_shader.n646[1] ));
 sg13g2_nor2_1 _3294_ (.A(\videogen.fancy_shader.video_y[1] ),
    .B(\videogen.fancy_shader.n646[1] ),
    .Y(_0986_));
 sg13g2_xor2_1 _3295_ (.B(\videogen.fancy_shader.n646[1] ),
    .A(\videogen.fancy_shader.video_y[1] ),
    .X(_0987_));
 sg13g2_nand2_1 _3296_ (.Y(_0988_),
    .A(net608),
    .B(\videogen.fancy_shader.n646[0] ));
 sg13g2_xor2_1 _3297_ (.B(\videogen.fancy_shader.n646[0] ),
    .A(net608),
    .X(_0989_));
 sg13g2_nand2_2 _3298_ (.Y(_0990_),
    .A(_0987_),
    .B(_0989_));
 sg13g2_o21ai_1 _3299_ (.B1(_0985_),
    .Y(_0991_),
    .A1(_0986_),
    .A2(_0988_));
 sg13g2_and2_1 _3300_ (.A(\videogen.fancy_shader.video_y[2] ),
    .B(\videogen.fancy_shader.n646[2] ),
    .X(_0992_));
 sg13g2_xor2_1 _3301_ (.B(\videogen.fancy_shader.n646[2] ),
    .A(\videogen.fancy_shader.video_y[2] ),
    .X(_0993_));
 sg13g2_xnor2_1 _3302_ (.Y(_0994_),
    .A(_0991_),
    .B(_0993_));
 sg13g2_nor2_2 _3303_ (.A(_0990_),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_nor2b_2 _3304_ (.A(_0942_),
    .B_N(_0995_),
    .Y(_0996_));
 sg13g2_nor3_1 _3305_ (.A(net750),
    .B(_0984_),
    .C(_0996_),
    .Y(_0348_));
 sg13g2_xnor2_1 _3306_ (.Y(_0997_),
    .A(\videogen.fancy_shader.n646[3] ),
    .B(_0996_));
 sg13g2_nor2_1 _3307_ (.A(net750),
    .B(_0997_),
    .Y(_0349_));
 sg13g2_nand2_1 _3308_ (.Y(_0998_),
    .A(\videogen.fancy_shader.n646[4] ),
    .B(\videogen.fancy_shader.video_x[4] ));
 sg13g2_xnor2_1 _3309_ (.Y(_0999_),
    .A(\videogen.fancy_shader.n646[4] ),
    .B(\videogen.fancy_shader.video_x[4] ));
 sg13g2_nor2_1 _3310_ (.A(\videogen.fancy_shader.n646[3] ),
    .B(\videogen.fancy_shader.video_x[3] ),
    .Y(_1000_));
 sg13g2_and2_1 _3311_ (.A(\videogen.fancy_shader.n646[2] ),
    .B(\videogen.fancy_shader.video_x[2] ),
    .X(_1001_));
 sg13g2_xor2_1 _3312_ (.B(\videogen.fancy_shader.video_x[2] ),
    .A(\videogen.fancy_shader.n646[2] ),
    .X(_1002_));
 sg13g2_nand2_1 _3313_ (.Y(_1003_),
    .A(\videogen.fancy_shader.n646[1] ),
    .B(\videogen.fancy_shader.video_x[1] ));
 sg13g2_nand2_1 _3314_ (.Y(_1004_),
    .A(\videogen.fancy_shader.n646[0] ),
    .B(\videogen.fancy_shader.video_x[0] ));
 sg13g2_xnor2_1 _3315_ (.Y(_1005_),
    .A(\videogen.fancy_shader.n646[1] ),
    .B(\videogen.fancy_shader.video_x[1] ));
 sg13g2_o21ai_1 _3316_ (.B1(_1003_),
    .Y(_1006_),
    .A1(_1004_),
    .A2(_1005_));
 sg13g2_a221oi_1 _3317_ (.B2(_1006_),
    .C1(_1001_),
    .B1(_1002_),
    .A1(\videogen.fancy_shader.n646[3] ),
    .Y(_1007_),
    .A2(\videogen.fancy_shader.video_x[3] ));
 sg13g2_or2_1 _3318_ (.X(_1008_),
    .B(_1007_),
    .A(_1000_));
 sg13g2_xnor2_1 _3319_ (.Y(_1009_),
    .A(_0999_),
    .B(_1008_));
 sg13g2_xnor2_1 _3320_ (.Y(_1010_),
    .A(\videogen.fancy_shader.n646[0] ),
    .B(\videogen.fancy_shader.video_x[0] ));
 sg13g2_nor2_2 _3321_ (.A(_1005_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_xor2_1 _3322_ (.B(_1006_),
    .A(_1002_),
    .X(_1012_));
 sg13g2_and2_1 _3323_ (.A(_1011_),
    .B(_1012_),
    .X(_1013_));
 sg13g2_xnor2_1 _3324_ (.Y(_1014_),
    .A(\videogen.fancy_shader.n646[3] ),
    .B(\videogen.fancy_shader.video_x[3] ));
 sg13g2_a21oi_1 _3325_ (.A1(_1002_),
    .A2(_1006_),
    .Y(_1015_),
    .B1(_1001_));
 sg13g2_xnor2_1 _3326_ (.Y(_1016_),
    .A(_1014_),
    .B(_1015_));
 sg13g2_nor2b_1 _3327_ (.A(_1016_),
    .B_N(_1013_),
    .Y(_1017_));
 sg13g2_nor2b_2 _3328_ (.A(_1009_),
    .B_N(_1017_),
    .Y(_1018_));
 sg13g2_nor2b_2 _3329_ (.A(_0942_),
    .B_N(_1018_),
    .Y(_1019_));
 sg13g2_a21oi_1 _3330_ (.A1(\videogen.fancy_shader.n646[3] ),
    .A2(_0996_),
    .Y(_1020_),
    .B1(\videogen.fancy_shader.n646[4] ));
 sg13g2_nor3_1 _3331_ (.A(net750),
    .B(_1019_),
    .C(_1020_),
    .Y(_0350_));
 sg13g2_xnor2_1 _3332_ (.Y(_1021_),
    .A(\videogen.fancy_shader.n646[5] ),
    .B(_1019_));
 sg13g2_nor2_1 _3333_ (.A(net745),
    .B(_1021_),
    .Y(_0351_));
 sg13g2_a21oi_1 _3334_ (.A1(\videogen.fancy_shader.n646[5] ),
    .A2(_1019_),
    .Y(_1022_),
    .B1(\videogen.fancy_shader.n646[6] ));
 sg13g2_nand3_1 _3335_ (.B(\videogen.fancy_shader.n646[5] ),
    .C(_1019_),
    .A(\videogen.fancy_shader.n646[6] ),
    .Y(_1023_));
 sg13g2_nand2_1 _3336_ (.Y(_1024_),
    .A(net795),
    .B(_1023_));
 sg13g2_nor2_1 _3337_ (.A(_1022_),
    .B(_1024_),
    .Y(_0352_));
 sg13g2_and2_1 _3338_ (.A(_0642_),
    .B(_1023_),
    .X(_1025_));
 sg13g2_nor2_1 _3339_ (.A(_0642_),
    .B(_1023_),
    .Y(_1026_));
 sg13g2_nor3_1 _3340_ (.A(net745),
    .B(_1025_),
    .C(_1026_),
    .Y(_0353_));
 sg13g2_or2_1 _3341_ (.X(_1027_),
    .B(_1026_),
    .A(net609));
 sg13g2_nand2_1 _3342_ (.Y(_1028_),
    .A(\videogen.fancy_shader.n646[8] ),
    .B(_1026_));
 sg13g2_and3_1 _3343_ (.X(_0354_),
    .A(net795),
    .B(_1027_),
    .C(_1028_));
 sg13g2_o21ai_1 _3344_ (.B1(net795),
    .Y(_1029_),
    .A1(_0641_),
    .A2(_1028_));
 sg13g2_a21oi_1 _3345_ (.A1(_0641_),
    .A2(_1028_),
    .Y(_0355_),
    .B1(_1029_));
 sg13g2_and2_1 _3346_ (.A(net608),
    .B(_0922_),
    .X(_1030_));
 sg13g2_o21ai_1 _3347_ (.B1(net797),
    .Y(_1031_),
    .A1(net608),
    .A2(_0922_));
 sg13g2_nor2_1 _3348_ (.A(_1030_),
    .B(_1031_),
    .Y(_0356_));
 sg13g2_and2_1 _3349_ (.A(\videogen.fancy_shader.video_y[1] ),
    .B(_1030_),
    .X(_1032_));
 sg13g2_nand2b_1 _3350_ (.Y(_1033_),
    .B(_0922_),
    .A_N(_0831_));
 sg13g2_o21ai_1 _3351_ (.B1(net798),
    .Y(_1034_),
    .A1(\videogen.fancy_shader.video_y[1] ),
    .A2(_1030_));
 sg13g2_nor2_1 _3352_ (.A(_1032_),
    .B(_1034_),
    .Y(_0357_));
 sg13g2_nor4_1 _3353_ (.A(\videogen.fancy_shader.video_y[7] ),
    .B(\videogen.fancy_shader.video_y[6] ),
    .C(\videogen.fancy_shader.video_y[5] ),
    .D(\videogen.fancy_shader.video_y[4] ),
    .Y(_1035_));
 sg13g2_nor4_1 _3354_ (.A(_0637_),
    .B(\videogen.fancy_shader.video_y[8] ),
    .C(_0831_),
    .D(_0935_),
    .Y(_1036_));
 sg13g2_nand3_1 _3355_ (.B(_1035_),
    .C(_1036_),
    .A(_0922_),
    .Y(_1037_));
 sg13g2_nand2_1 _3356_ (.Y(_1038_),
    .A(net797),
    .B(_1037_));
 sg13g2_xnor2_1 _3357_ (.Y(_1039_),
    .A(_0640_),
    .B(_1033_));
 sg13g2_nor2_1 _3358_ (.A(_1038_),
    .B(_1039_),
    .Y(_0358_));
 sg13g2_a22oi_1 _3359_ (.Y(_1040_),
    .B1(_1037_),
    .B2(\videogen.fancy_shader.video_y[3] ),
    .A2(_1032_),
    .A1(\videogen.fancy_shader.video_y[2] ));
 sg13g2_nor2_1 _3360_ (.A(_0829_),
    .B(_1033_),
    .Y(_1041_));
 sg13g2_nor3_1 _3361_ (.A(net750),
    .B(_1040_),
    .C(_1041_),
    .Y(_0359_));
 sg13g2_nor2_1 _3362_ (.A(\videogen.fancy_shader.video_y[4] ),
    .B(_1041_),
    .Y(_1042_));
 sg13g2_nand3_1 _3363_ (.B(_0834_),
    .C(_0922_),
    .A(\videogen.fancy_shader.video_y[4] ),
    .Y(_1043_));
 sg13g2_and2_1 _3364_ (.A(\videogen.fancy_shader.video_y[4] ),
    .B(_1041_),
    .X(_1044_));
 sg13g2_nor3_1 _3365_ (.A(net745),
    .B(_1042_),
    .C(_1044_),
    .Y(_0360_));
 sg13g2_nor2_1 _3366_ (.A(\videogen.fancy_shader.video_y[5] ),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_and2_1 _3367_ (.A(\videogen.fancy_shader.video_y[5] ),
    .B(_1044_),
    .X(_1046_));
 sg13g2_nor3_1 _3368_ (.A(net745),
    .B(_1045_),
    .C(_1046_),
    .Y(_0361_));
 sg13g2_xnor2_1 _3369_ (.Y(_1047_),
    .A(\videogen.fancy_shader.video_y[6] ),
    .B(_1046_));
 sg13g2_nor2_1 _3370_ (.A(net746),
    .B(_1047_),
    .Y(_0362_));
 sg13g2_a21oi_1 _3371_ (.A1(\videogen.fancy_shader.video_y[6] ),
    .A2(_1046_),
    .Y(_1048_),
    .B1(\videogen.fancy_shader.video_y[7] ));
 sg13g2_nor2_1 _3372_ (.A(_0673_),
    .B(_1043_),
    .Y(_1049_));
 sg13g2_nor3_1 _3373_ (.A(net745),
    .B(_1048_),
    .C(_1049_),
    .Y(_0363_));
 sg13g2_nor2_1 _3374_ (.A(\videogen.fancy_shader.video_y[8] ),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_nor3_1 _3375_ (.A(_0638_),
    .B(_0673_),
    .C(_1043_),
    .Y(_1051_));
 sg13g2_nor3_1 _3376_ (.A(net745),
    .B(_1050_),
    .C(_1051_),
    .Y(_0364_));
 sg13g2_xnor2_1 _3377_ (.Y(_1052_),
    .A(\videogen.fancy_shader.video_y[9] ),
    .B(_1051_));
 sg13g2_nor2_1 _3378_ (.A(_1038_),
    .B(_1052_),
    .Y(_0365_));
 sg13g2_nor2_1 _3379_ (.A(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .B(net746),
    .Y(_0366_));
 sg13g2_o21ai_1 _3380_ (.B1(net796),
    .Y(_1053_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ));
 sg13g2_a21oi_1 _3381_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .Y(_0367_),
    .B1(_1053_));
 sg13g2_a21oi_1 _3382_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .Y(_1054_),
    .B1(\videogen.test_lut_thingy.gol_counter_reg[2] ));
 sg13g2_and3_1 _3383_ (.X(_1055_),
    .A(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .B(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .C(\videogen.test_lut_thingy.gol_counter_reg[2] ));
 sg13g2_nor3_1 _3384_ (.A(net751),
    .B(_1054_),
    .C(_1055_),
    .Y(_0368_));
 sg13g2_o21ai_1 _3385_ (.B1(net795),
    .Y(_1056_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A2(_1055_));
 sg13g2_a21oi_1 _3386_ (.A1(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A2(_1055_),
    .Y(_0369_),
    .B1(_1056_));
 sg13g2_nand4_1 _3387_ (.B(\videogen.fancy_shader.video_x[6] ),
    .C(\videogen.fancy_shader.video_x[5] ),
    .A(\videogen.fancy_shader.video_x[7] ),
    .Y(_1057_),
    .D(_0926_));
 sg13g2_a21oi_1 _3388_ (.A1(_0678_),
    .A2(_0813_),
    .Y(_1058_),
    .B1(_0805_));
 sg13g2_a21oi_1 _3389_ (.A1(_1057_),
    .A2(_1058_),
    .Y(_0370_),
    .B1(net745));
 sg13g2_xnor2_1 _3390_ (.Y(_1059_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_xor2_1 _3391_ (.B(_1005_),
    .A(_1004_),
    .X(_1060_));
 sg13g2_nand2_1 _3392_ (.Y(_1061_),
    .A(_1059_),
    .B(_1060_));
 sg13g2_or2_1 _3393_ (.X(_1062_),
    .B(_1060_),
    .A(_1059_));
 sg13g2_and2_1 _3394_ (.A(_1061_),
    .B(_1062_),
    .X(_1063_));
 sg13g2_inv_1 _3395_ (.Y(_1064_),
    .A(_1063_));
 sg13g2_xnor2_1 _3396_ (.Y(_1065_),
    .A(_0994_),
    .B(_1012_));
 sg13g2_inv_2 _3397_ (.Y(_1066_),
    .A(_1065_));
 sg13g2_nor2_1 _3398_ (.A(\videogen.fancy_shader.video_y[3] ),
    .B(\videogen.fancy_shader.n646[3] ),
    .Y(_1067_));
 sg13g2_a221oi_1 _3399_ (.B2(_0993_),
    .C1(_0992_),
    .B1(_0991_),
    .A1(\videogen.fancy_shader.video_y[3] ),
    .Y(_1068_),
    .A2(\videogen.fancy_shader.n646[3] ));
 sg13g2_nand2_1 _3400_ (.Y(_1069_),
    .A(\videogen.fancy_shader.video_y[4] ),
    .B(\videogen.fancy_shader.n646[4] ));
 sg13g2_xnor2_1 _3401_ (.Y(_1070_),
    .A(\videogen.fancy_shader.video_y[4] ),
    .B(\videogen.fancy_shader.n646[4] ));
 sg13g2_or3_1 _3402_ (.A(_1067_),
    .B(_1068_),
    .C(_1070_),
    .X(_1071_));
 sg13g2_o21ai_1 _3403_ (.B1(_1070_),
    .Y(_1072_),
    .A1(_1067_),
    .A2(_1068_));
 sg13g2_nand2_2 _3404_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_or2_1 _3405_ (.X(_1074_),
    .B(_1073_),
    .A(_1009_));
 sg13g2_nand2_1 _3406_ (.Y(_1075_),
    .A(_1009_),
    .B(_1073_));
 sg13g2_nand2_2 _3407_ (.Y(_1076_),
    .A(_1074_),
    .B(_1075_));
 sg13g2_and2_1 _3408_ (.A(_1074_),
    .B(_1075_),
    .X(_1077_));
 sg13g2_nor2_1 _3409_ (.A(\videogen.fancy_shader.n646[5] ),
    .B(\videogen.fancy_shader.video_x[5] ),
    .Y(_1078_));
 sg13g2_nand2_1 _3410_ (.Y(_1079_),
    .A(\videogen.fancy_shader.n646[5] ),
    .B(\videogen.fancy_shader.video_x[5] ));
 sg13g2_nand2b_1 _3411_ (.Y(_1080_),
    .B(_1079_),
    .A_N(_1078_));
 sg13g2_o21ai_1 _3412_ (.B1(_0998_),
    .Y(_1081_),
    .A1(_0999_),
    .A2(_1008_));
 sg13g2_xnor2_1 _3413_ (.Y(_1082_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_nor2_1 _3414_ (.A(\videogen.fancy_shader.video_y[5] ),
    .B(\videogen.fancy_shader.n646[5] ),
    .Y(_1083_));
 sg13g2_nand2_1 _3415_ (.Y(_1084_),
    .A(\videogen.fancy_shader.video_y[5] ),
    .B(\videogen.fancy_shader.n646[5] ));
 sg13g2_nand2b_1 _3416_ (.Y(_1085_),
    .B(_1084_),
    .A_N(_1083_));
 sg13g2_and3_1 _3417_ (.X(_1086_),
    .A(_1069_),
    .B(_1071_),
    .C(_1085_));
 sg13g2_a21oi_1 _3418_ (.A1(_1069_),
    .A2(_1071_),
    .Y(_1087_),
    .B1(_1085_));
 sg13g2_nor2_1 _3419_ (.A(_1086_),
    .B(_1087_),
    .Y(_1088_));
 sg13g2_xor2_1 _3420_ (.B(_1088_),
    .A(_1082_),
    .X(_1089_));
 sg13g2_inv_1 _3421_ (.Y(_1090_),
    .A(net544));
 sg13g2_and2_1 _3422_ (.A(\videogen.fancy_shader.video_y[8] ),
    .B(net609),
    .X(_1091_));
 sg13g2_nand2_1 _3423_ (.Y(_1092_),
    .A(\videogen.fancy_shader.video_y[8] ),
    .B(net609));
 sg13g2_or2_1 _3424_ (.X(_1093_),
    .B(_1085_),
    .A(_1070_));
 sg13g2_nor3_1 _3425_ (.A(_1067_),
    .B(_1068_),
    .C(_1093_),
    .Y(_1094_));
 sg13g2_a21oi_1 _3426_ (.A1(_1069_),
    .A2(_1084_),
    .Y(_1095_),
    .B1(_1083_));
 sg13g2_xor2_1 _3427_ (.B(\videogen.fancy_shader.n646[7] ),
    .A(\videogen.fancy_shader.video_y[7] ),
    .X(_1096_));
 sg13g2_xnor2_1 _3428_ (.Y(_1097_),
    .A(\videogen.fancy_shader.video_y[7] ),
    .B(\videogen.fancy_shader.n646[7] ));
 sg13g2_nand2_2 _3429_ (.Y(_1098_),
    .A(\videogen.fancy_shader.video_y[6] ),
    .B(\videogen.fancy_shader.n646[6] ));
 sg13g2_xor2_1 _3430_ (.B(\videogen.fancy_shader.n646[6] ),
    .A(\videogen.fancy_shader.video_y[6] ),
    .X(_1099_));
 sg13g2_and2_1 _3431_ (.A(_1096_),
    .B(_1099_),
    .X(_1100_));
 sg13g2_o21ai_1 _3432_ (.B1(_1100_),
    .Y(_1101_),
    .A1(_1094_),
    .A2(_1095_));
 sg13g2_a21oi_1 _3433_ (.A1(_0639_),
    .A2(_0642_),
    .Y(_1102_),
    .B1(_1098_));
 sg13g2_a21oi_2 _3434_ (.B1(_1102_),
    .Y(_1103_),
    .A2(\videogen.fancy_shader.n646[7] ),
    .A1(\videogen.fancy_shader.video_y[7] ));
 sg13g2_xor2_1 _3435_ (.B(net609),
    .A(\videogen.fancy_shader.video_y[8] ),
    .X(_1104_));
 sg13g2_xnor2_1 _3436_ (.Y(_1105_),
    .A(\videogen.fancy_shader.video_y[8] ),
    .B(net609));
 sg13g2_a21oi_1 _3437_ (.A1(_1101_),
    .A2(_1103_),
    .Y(_1106_),
    .B1(_1105_));
 sg13g2_a21o_1 _3438_ (.A2(_1103_),
    .A1(_1101_),
    .B1(_1105_),
    .X(_1107_));
 sg13g2_xnor2_1 _3439_ (.Y(_1108_),
    .A(\videogen.fancy_shader.video_y[9] ),
    .B(\videogen.fancy_shader.n646[9] ));
 sg13g2_xor2_1 _3440_ (.B(\videogen.fancy_shader.n646[9] ),
    .A(\videogen.fancy_shader.video_y[9] ),
    .X(_1109_));
 sg13g2_nand3_1 _3441_ (.B(_1107_),
    .C(_1109_),
    .A(_1092_),
    .Y(_1110_));
 sg13g2_o21ai_1 _3442_ (.B1(_1108_),
    .Y(_1111_),
    .A1(_1091_),
    .A2(_1106_));
 sg13g2_nand3_1 _3443_ (.B(_1107_),
    .C(_1108_),
    .A(_1092_),
    .Y(_1112_));
 sg13g2_o21ai_1 _3444_ (.B1(_1109_),
    .Y(_1113_),
    .A1(_1091_),
    .A2(_1106_));
 sg13g2_and2_1 _3445_ (.A(net609),
    .B(\videogen.fancy_shader.video_x[8] ),
    .X(_1114_));
 sg13g2_nand2_1 _3446_ (.Y(_1115_),
    .A(net609),
    .B(\videogen.fancy_shader.video_x[8] ));
 sg13g2_nor4_1 _3447_ (.A(_0999_),
    .B(_1000_),
    .C(_1007_),
    .D(_1080_),
    .Y(_1116_));
 sg13g2_a21oi_1 _3448_ (.A1(_0998_),
    .A2(_1079_),
    .Y(_1117_),
    .B1(_1078_));
 sg13g2_xnor2_1 _3449_ (.Y(_1118_),
    .A(\videogen.fancy_shader.n646[7] ),
    .B(net629));
 sg13g2_nand2_1 _3450_ (.Y(_1119_),
    .A(\videogen.fancy_shader.n646[6] ),
    .B(\videogen.fancy_shader.video_x[6] ));
 sg13g2_xor2_1 _3451_ (.B(\videogen.fancy_shader.video_x[6] ),
    .A(\videogen.fancy_shader.n646[6] ),
    .X(_1120_));
 sg13g2_nor2b_1 _3452_ (.A(_1118_),
    .B_N(_1120_),
    .Y(_1121_));
 sg13g2_o21ai_1 _3453_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_a21oi_1 _3454_ (.A1(_0642_),
    .A2(_0651_),
    .Y(_1123_),
    .B1(_1119_));
 sg13g2_a21oi_1 _3455_ (.A1(\videogen.fancy_shader.n646[7] ),
    .A2(net629),
    .Y(_1124_),
    .B1(_1123_));
 sg13g2_xnor2_1 _3456_ (.Y(_1125_),
    .A(net609),
    .B(\videogen.fancy_shader.video_x[8] ));
 sg13g2_a21oi_1 _3457_ (.A1(_1122_),
    .A2(_1124_),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_a21o_2 _3458_ (.A2(_1124_),
    .A1(_1122_),
    .B1(_1125_),
    .X(_1127_));
 sg13g2_xor2_1 _3459_ (.B(\videogen.fancy_shader.video_x[9] ),
    .A(\videogen.fancy_shader.n646[9] ),
    .X(_1128_));
 sg13g2_xnor2_1 _3460_ (.Y(_1129_),
    .A(\videogen.fancy_shader.n646[9] ),
    .B(\videogen.fancy_shader.video_x[9] ));
 sg13g2_nand3_1 _3461_ (.B(_1127_),
    .C(_1129_),
    .A(_1115_),
    .Y(_1130_));
 sg13g2_o21ai_1 _3462_ (.B1(_1128_),
    .Y(_1131_),
    .A1(_1114_),
    .A2(_1126_));
 sg13g2_o21ai_1 _3463_ (.B1(_1129_),
    .Y(_1132_),
    .A1(_1114_),
    .A2(_1126_));
 sg13g2_nand3_1 _3464_ (.B(_1127_),
    .C(_1128_),
    .A(_1115_),
    .Y(_1133_));
 sg13g2_a22oi_1 _3465_ (.Y(_1134_),
    .B1(_1130_),
    .B2(_1131_),
    .A2(_1113_),
    .A1(_1112_));
 sg13g2_nand4_1 _3466_ (.B(_1111_),
    .C(_1132_),
    .A(_1110_),
    .Y(_1135_),
    .D(_1133_));
 sg13g2_a22oi_1 _3467_ (.Y(_1136_),
    .B1(_1132_),
    .B2(_1133_),
    .A2(_1111_),
    .A1(_1110_));
 sg13g2_nand4_1 _3468_ (.B(_1113_),
    .C(_1130_),
    .A(_1112_),
    .Y(_1137_),
    .D(_1131_));
 sg13g2_nand2_1 _3469_ (.Y(_1138_),
    .A(_1135_),
    .B(_1137_));
 sg13g2_nor2_2 _3470_ (.A(_1134_),
    .B(_1136_),
    .Y(_1139_));
 sg13g2_o21ai_1 _3471_ (.B1(_1120_),
    .Y(_1140_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_or3_1 _3472_ (.A(_1116_),
    .B(_1117_),
    .C(_1120_),
    .X(_1141_));
 sg13g2_and2_1 _3473_ (.A(_1140_),
    .B(_1141_),
    .X(_1142_));
 sg13g2_o21ai_1 _3474_ (.B1(_1099_),
    .Y(_1143_),
    .A1(_1094_),
    .A2(_1095_));
 sg13g2_or3_1 _3475_ (.A(_1094_),
    .B(_1095_),
    .C(_1099_),
    .X(_1144_));
 sg13g2_and2_1 _3476_ (.A(_1143_),
    .B(_1144_),
    .X(_1145_));
 sg13g2_xor2_1 _3477_ (.B(_1145_),
    .A(_1142_),
    .X(_1146_));
 sg13g2_xnor2_1 _3478_ (.Y(_1147_),
    .A(_1142_),
    .B(_1145_));
 sg13g2_a21oi_2 _3479_ (.B1(_1147_),
    .Y(_1148_),
    .A2(_1137_),
    .A1(_1135_));
 sg13g2_nor3_1 _3480_ (.A(_1134_),
    .B(_1136_),
    .C(_1146_),
    .Y(_1149_));
 sg13g2_nand3_1 _3481_ (.B(_1119_),
    .C(_1140_),
    .A(_1118_),
    .Y(_1150_));
 sg13g2_a21o_1 _3482_ (.A2(_1140_),
    .A1(_1119_),
    .B1(_1118_),
    .X(_1151_));
 sg13g2_nand3_1 _3483_ (.B(_1098_),
    .C(_1143_),
    .A(_1096_),
    .Y(_1152_));
 sg13g2_a21o_1 _3484_ (.A2(_1143_),
    .A1(_1098_),
    .B1(_1096_),
    .X(_1153_));
 sg13g2_nand3_1 _3485_ (.B(_1098_),
    .C(_1143_),
    .A(_1097_),
    .Y(_1154_));
 sg13g2_a21o_1 _3486_ (.A2(_1143_),
    .A1(_1098_),
    .B1(_1097_),
    .X(_1155_));
 sg13g2_a22oi_1 _3487_ (.Y(_1156_),
    .B1(_1152_),
    .B2(_1153_),
    .A2(_1151_),
    .A1(_1150_));
 sg13g2_and4_1 _3488_ (.A(_1150_),
    .B(_1151_),
    .C(_1152_),
    .D(_1153_),
    .X(_1157_));
 sg13g2_nor2_2 _3489_ (.A(_1156_),
    .B(_1157_),
    .Y(_1158_));
 sg13g2_nand3_1 _3490_ (.B(_1124_),
    .C(_1125_),
    .A(_1122_),
    .Y(_1159_));
 sg13g2_nand2_1 _3491_ (.Y(_1160_),
    .A(_1127_),
    .B(_1159_));
 sg13g2_nand3_1 _3492_ (.B(_1103_),
    .C(_1104_),
    .A(_1101_),
    .Y(_1161_));
 sg13g2_a21o_2 _3493_ (.A2(_1103_),
    .A1(_1101_),
    .B1(_1104_),
    .X(_1162_));
 sg13g2_nand2_1 _3494_ (.Y(_1163_),
    .A(_1161_),
    .B(_1162_));
 sg13g2_a22oi_1 _3495_ (.Y(_1164_),
    .B1(_1161_),
    .B2(_1162_),
    .A2(_1159_),
    .A1(_1127_));
 sg13g2_and4_1 _3496_ (.A(_1127_),
    .B(_1159_),
    .C(_1161_),
    .D(_1162_),
    .X(_1165_));
 sg13g2_or2_1 _3497_ (.X(_1166_),
    .B(_1165_),
    .A(_1164_));
 sg13g2_nor2_1 _3498_ (.A(_1164_),
    .B(_1165_),
    .Y(_1167_));
 sg13g2_nor4_1 _3499_ (.A(_1156_),
    .B(_1157_),
    .C(_1164_),
    .D(_1165_),
    .Y(_1168_));
 sg13g2_nor4_1 _3500_ (.A(_1134_),
    .B(_1136_),
    .C(_1146_),
    .D(_1168_),
    .Y(_1169_));
 sg13g2_or2_1 _3501_ (.X(_1170_),
    .B(_1169_),
    .A(_1148_));
 sg13g2_nand2_1 _3502_ (.Y(_1171_),
    .A(_1090_),
    .B(_1158_));
 sg13g2_or3_1 _3503_ (.A(_1148_),
    .B(_1169_),
    .C(_1171_),
    .X(_1172_));
 sg13g2_nor2_2 _3504_ (.A(_1158_),
    .B(_1167_),
    .Y(_1173_));
 sg13g2_a21oi_1 _3505_ (.A1(_1149_),
    .A2(_1158_),
    .Y(_1174_),
    .B1(_1167_));
 sg13g2_and2_1 _3506_ (.A(_1149_),
    .B(_1168_),
    .X(_1175_));
 sg13g2_a21oi_1 _3507_ (.A1(_1172_),
    .A2(_1174_),
    .Y(_1176_),
    .B1(_1175_));
 sg13g2_nor2_1 _3508_ (.A(net544),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_xnor2_1 _3509_ (.Y(_1178_),
    .A(net544),
    .B(_1176_));
 sg13g2_nor3_1 _3510_ (.A(_1077_),
    .B(_1170_),
    .C(_1178_),
    .Y(_1179_));
 sg13g2_nor3_1 _3511_ (.A(net544),
    .B(_1170_),
    .C(_1176_),
    .Y(_1180_));
 sg13g2_or3_1 _3512_ (.A(_1149_),
    .B(_1158_),
    .C(_1180_),
    .X(_1181_));
 sg13g2_o21ai_1 _3513_ (.B1(_1158_),
    .Y(_1182_),
    .A1(_1169_),
    .A2(_1180_));
 sg13g2_and2_1 _3514_ (.A(_1181_),
    .B(_1182_),
    .X(_1183_));
 sg13g2_a21o_1 _3515_ (.A2(_1182_),
    .A1(_1181_),
    .B1(_1179_),
    .X(_1184_));
 sg13g2_nor2b_1 _3516_ (.A(_1172_),
    .B_N(_1174_),
    .Y(_1185_));
 sg13g2_a21oi_2 _3517_ (.B1(_1185_),
    .Y(_1186_),
    .A2(_1175_),
    .A1(net544));
 sg13g2_a21o_1 _3518_ (.A2(_1186_),
    .A1(_1184_),
    .B1(_1077_),
    .X(_1187_));
 sg13g2_nand3_1 _3519_ (.B(_1184_),
    .C(_1186_),
    .A(_1077_),
    .Y(_1188_));
 sg13g2_nand2_1 _3520_ (.Y(_1189_),
    .A(_1187_),
    .B(_1188_));
 sg13g2_xor2_1 _3521_ (.B(\videogen.fancy_shader.n646[3] ),
    .A(\videogen.fancy_shader.video_y[3] ),
    .X(_1190_));
 sg13g2_a21oi_1 _3522_ (.A1(_0991_),
    .A2(_0993_),
    .Y(_1191_),
    .B1(_0992_));
 sg13g2_xnor2_1 _3523_ (.Y(_1192_),
    .A(_1190_),
    .B(_1191_));
 sg13g2_nand2b_1 _3524_ (.Y(_1193_),
    .B(_1192_),
    .A_N(_1016_));
 sg13g2_nand2b_1 _3525_ (.Y(_1194_),
    .B(_1016_),
    .A_N(_1192_));
 sg13g2_and2_1 _3526_ (.A(_1193_),
    .B(_1194_),
    .X(_1195_));
 sg13g2_nand2_1 _3527_ (.Y(_1196_),
    .A(_1193_),
    .B(_1194_));
 sg13g2_nor2_1 _3528_ (.A(_1178_),
    .B(_1195_),
    .Y(_1197_));
 sg13g2_nand3_1 _3529_ (.B(_1188_),
    .C(_1197_),
    .A(_1187_),
    .Y(_1198_));
 sg13g2_o21ai_1 _3530_ (.B1(_1183_),
    .Y(_1199_),
    .A1(_1179_),
    .A2(_1186_));
 sg13g2_and2_1 _3531_ (.A(_1184_),
    .B(_1199_),
    .X(_1200_));
 sg13g2_inv_1 _3532_ (.Y(_1201_),
    .A(_1200_));
 sg13g2_a221oi_1 _3533_ (.B2(_1186_),
    .C1(_1178_),
    .B1(_1184_),
    .A1(_1074_),
    .Y(_1202_),
    .A2(_1075_));
 sg13g2_or3_1 _3534_ (.A(_1170_),
    .B(_1177_),
    .C(_1202_),
    .X(_1203_));
 sg13g2_o21ai_1 _3535_ (.B1(_1170_),
    .Y(_1204_),
    .A1(_1177_),
    .A2(_1202_));
 sg13g2_nand2_1 _3536_ (.Y(_1205_),
    .A(_1203_),
    .B(_1204_));
 sg13g2_nand3_1 _3537_ (.B(_1203_),
    .C(_1204_),
    .A(_1198_),
    .Y(_1206_));
 sg13g2_nand2b_1 _3538_ (.Y(_1207_),
    .B(_1200_),
    .A_N(_1198_));
 sg13g2_a21o_1 _3539_ (.A2(_1206_),
    .A1(_1201_),
    .B1(_1195_),
    .X(_1208_));
 sg13g2_a221oi_1 _3540_ (.B2(_1206_),
    .C1(_1189_),
    .B1(_1201_),
    .A1(_1193_),
    .Y(_1209_),
    .A2(_1194_));
 sg13g2_xor2_1 _3541_ (.B(_1187_),
    .A(_1178_),
    .X(_1210_));
 sg13g2_o21ai_1 _3542_ (.B1(_1207_),
    .Y(_1211_),
    .A1(_1209_),
    .A2(_1210_));
 sg13g2_nand3_1 _3543_ (.B(_1201_),
    .C(_1205_),
    .A(_1195_),
    .Y(_1212_));
 sg13g2_and2_1 _3544_ (.A(_1208_),
    .B(_1212_),
    .X(_1213_));
 sg13g2_nor2_1 _3545_ (.A(_1065_),
    .B(_1189_),
    .Y(_1214_));
 sg13g2_nand3_1 _3546_ (.B(_1212_),
    .C(_1214_),
    .A(_1208_),
    .Y(_1215_));
 sg13g2_nand2_1 _3547_ (.Y(_1216_),
    .A(_1198_),
    .B(_1200_));
 sg13g2_o21ai_1 _3548_ (.B1(_1216_),
    .Y(_1217_),
    .A1(_1198_),
    .A2(_1205_));
 sg13g2_a21oi_1 _3549_ (.A1(_1211_),
    .A2(_1215_),
    .Y(_1218_),
    .B1(_1217_));
 sg13g2_nor2_1 _3550_ (.A(_1065_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_xnor2_1 _3551_ (.Y(_1220_),
    .A(_1065_),
    .B(_1218_));
 sg13g2_nand2_1 _3552_ (.Y(_1221_),
    .A(_1064_),
    .B(_1213_));
 sg13g2_or2_1 _3553_ (.X(_1222_),
    .B(_1221_),
    .A(_1220_));
 sg13g2_nand3b_1 _3554_ (.B(_1213_),
    .C(_1066_),
    .Y(_1223_),
    .A_N(_1218_));
 sg13g2_a21oi_1 _3555_ (.A1(_1208_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(_1189_));
 sg13g2_and3_1 _3556_ (.X(_1225_),
    .A(_1189_),
    .B(_1208_),
    .C(_1223_));
 sg13g2_or2_1 _3557_ (.X(_1226_),
    .B(_1225_),
    .A(_1224_));
 sg13g2_o21ai_1 _3558_ (.B1(_1222_),
    .Y(_1227_),
    .A1(_1224_),
    .A2(_1225_));
 sg13g2_a21oi_1 _3559_ (.A1(_1215_),
    .A2(_1217_),
    .Y(_1228_),
    .B1(_1211_));
 sg13g2_a21oi_1 _3560_ (.A1(_1211_),
    .A2(_1215_),
    .Y(_1229_),
    .B1(_1228_));
 sg13g2_a21o_1 _3561_ (.A2(_1215_),
    .A1(_1211_),
    .B1(_1228_),
    .X(_1230_));
 sg13g2_and2_1 _3562_ (.A(_1227_),
    .B(_1230_),
    .X(_1231_));
 sg13g2_xnor2_1 _3563_ (.Y(_1232_),
    .A(_1063_),
    .B(_1231_));
 sg13g2_or2_1 _3564_ (.X(_1233_),
    .B(\videogen.fancy_shader.video_x[0] ),
    .A(net608));
 sg13g2_nand2_1 _3565_ (.Y(_1234_),
    .A(\videogen.fancy_shader.video_y[0] ),
    .B(\videogen.fancy_shader.video_x[0] ));
 sg13g2_nand2_2 _3566_ (.Y(_1235_),
    .A(_1233_),
    .B(_1234_));
 sg13g2_and2_1 _3567_ (.A(_1233_),
    .B(_1234_),
    .X(_1236_));
 sg13g2_nor2b_1 _3568_ (.A(_1222_),
    .B_N(_1226_),
    .Y(_1237_));
 sg13g2_a21oi_1 _3569_ (.A1(_1222_),
    .A2(_1229_),
    .Y(_1238_),
    .B1(_1237_));
 sg13g2_a221oi_1 _3570_ (.B2(_1230_),
    .C1(_1220_),
    .B1(_1227_),
    .A1(_1061_),
    .Y(_1239_),
    .A2(_1062_));
 sg13g2_or3_1 _3571_ (.A(_1213_),
    .B(_1219_),
    .C(_1239_),
    .X(_1240_));
 sg13g2_o21ai_1 _3572_ (.B1(_1213_),
    .Y(_1241_),
    .A1(_1219_),
    .A2(_1239_));
 sg13g2_and3_1 _3573_ (.X(_1242_),
    .A(_1238_),
    .B(_1240_),
    .C(_1241_));
 sg13g2_o21ai_1 _3574_ (.B1(_1232_),
    .Y(_1243_),
    .A1(_1236_),
    .A2(_1242_));
 sg13g2_a221oi_1 _3575_ (.B2(_1241_),
    .C1(_1232_),
    .B1(_1240_),
    .A1(_1233_),
    .Y(_1244_),
    .A2(_1234_));
 sg13g2_o21ai_1 _3576_ (.B1(_1220_),
    .Y(_1245_),
    .A1(_1063_),
    .A2(_1231_));
 sg13g2_nor2_1 _3577_ (.A(_1138_),
    .B(_1173_),
    .Y(_1246_));
 sg13g2_mux2_1 _3578_ (.A0(_1139_),
    .A1(_1148_),
    .S(_1173_),
    .X(_1247_));
 sg13g2_and2_1 _3579_ (.A(_1146_),
    .B(_1247_),
    .X(_1248_));
 sg13g2_nor2_1 _3580_ (.A(_1146_),
    .B(_1246_),
    .Y(_1249_));
 sg13g2_nor2_2 _3581_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_a21oi_1 _3582_ (.A1(_1139_),
    .A2(_1166_),
    .Y(_1251_),
    .B1(_1158_));
 sg13g2_nand2_1 _3583_ (.Y(_1252_),
    .A(net544),
    .B(_1251_));
 sg13g2_nor3_1 _3584_ (.A(_1248_),
    .B(_1249_),
    .C(_1252_),
    .Y(_1253_));
 sg13g2_nand3_1 _3585_ (.B(_1247_),
    .C(_1251_),
    .A(_1146_),
    .Y(_1254_));
 sg13g2_xnor2_1 _3586_ (.Y(_1255_),
    .A(_1248_),
    .B(_1251_));
 sg13g2_o21ai_1 _3587_ (.B1(_1166_),
    .Y(_1256_),
    .A1(_1138_),
    .A2(_1158_));
 sg13g2_a22oi_1 _3588_ (.Y(_1257_),
    .B1(_1254_),
    .B2(_1256_),
    .A2(_1173_),
    .A1(_1148_));
 sg13g2_a221oi_1 _3589_ (.B2(_1256_),
    .C1(_1090_),
    .B1(_1254_),
    .A1(_1148_),
    .Y(_1258_),
    .A2(_1173_));
 sg13g2_or2_1 _3590_ (.X(_1259_),
    .B(_1258_),
    .A(_1253_));
 sg13g2_o21ai_1 _3591_ (.B1(_1250_),
    .Y(_1260_),
    .A1(_1253_),
    .A2(_1258_));
 sg13g2_a21oi_1 _3592_ (.A1(_1255_),
    .A2(_1260_),
    .Y(_1261_),
    .B1(_1253_));
 sg13g2_nor2_1 _3593_ (.A(net544),
    .B(_1257_),
    .Y(_1262_));
 sg13g2_or2_1 _3594_ (.X(_1263_),
    .B(_1262_),
    .A(_1259_));
 sg13g2_nor3_1 _3595_ (.A(_1076_),
    .B(_1259_),
    .C(_1262_),
    .Y(_1264_));
 sg13g2_a21oi_1 _3596_ (.A1(_1250_),
    .A2(_1264_),
    .Y(_1265_),
    .B1(_1261_));
 sg13g2_nor2_1 _3597_ (.A(_1076_),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_xnor2_1 _3598_ (.Y(_1267_),
    .A(_1076_),
    .B(_1265_));
 sg13g2_inv_1 _3599_ (.Y(_1268_),
    .A(_1267_));
 sg13g2_o21ai_1 _3600_ (.B1(_1264_),
    .Y(_1269_),
    .A1(_1250_),
    .A2(_1261_));
 sg13g2_o21ai_1 _3601_ (.B1(_1260_),
    .Y(_1270_),
    .A1(_1250_),
    .A2(_1258_));
 sg13g2_xnor2_1 _3602_ (.Y(_1271_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_o21ai_1 _3603_ (.B1(_1271_),
    .Y(_1272_),
    .A1(_1263_),
    .A2(_1267_));
 sg13g2_and2_1 _3604_ (.A(_1195_),
    .B(_1272_),
    .X(_1273_));
 sg13g2_and2_1 _3605_ (.A(_1196_),
    .B(_1271_),
    .X(_1274_));
 sg13g2_nor2_1 _3606_ (.A(_1273_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_nor3_1 _3607_ (.A(_1066_),
    .B(_1273_),
    .C(_1274_),
    .Y(_1276_));
 sg13g2_a21oi_1 _3608_ (.A1(_1268_),
    .A2(_1273_),
    .Y(_1277_),
    .B1(_1266_));
 sg13g2_xor2_1 _3609_ (.B(_1277_),
    .A(_1263_),
    .X(_1278_));
 sg13g2_a21o_1 _3610_ (.A2(_1276_),
    .A1(_1268_),
    .B1(_1278_),
    .X(_1279_));
 sg13g2_a21oi_1 _3611_ (.A1(_1276_),
    .A2(_1279_),
    .Y(_1280_),
    .B1(_1273_));
 sg13g2_xnor2_1 _3612_ (.Y(_1281_),
    .A(_1267_),
    .B(_1280_));
 sg13g2_xnor2_1 _3613_ (.Y(_1282_),
    .A(_1066_),
    .B(_1279_));
 sg13g2_nand2_1 _3614_ (.Y(_1283_),
    .A(_1275_),
    .B(_1282_));
 sg13g2_a21oi_1 _3615_ (.A1(_1281_),
    .A2(_1283_),
    .Y(_1284_),
    .B1(_1064_));
 sg13g2_and2_1 _3616_ (.A(_1064_),
    .B(_1281_),
    .X(_1285_));
 sg13g2_nand2_1 _3617_ (.Y(_1286_),
    .A(_1236_),
    .B(_1282_));
 sg13g2_nor3_1 _3618_ (.A(_1284_),
    .B(_1285_),
    .C(_1286_),
    .Y(_1287_));
 sg13g2_nor2_1 _3619_ (.A(_1235_),
    .B(_1275_),
    .Y(_1288_));
 sg13g2_nor2b_1 _3620_ (.A(_1288_),
    .B_N(_1282_),
    .Y(_1289_));
 sg13g2_a21o_1 _3621_ (.A2(_1278_),
    .A1(_1065_),
    .B1(_1275_),
    .X(_1290_));
 sg13g2_a21oi_1 _3622_ (.A1(_1276_),
    .A2(_1279_),
    .Y(_1291_),
    .B1(_1235_));
 sg13g2_a21oi_1 _3623_ (.A1(_1290_),
    .A2(_1291_),
    .Y(_1292_),
    .B1(_1282_));
 sg13g2_a22oi_1 _3624_ (.Y(_1293_),
    .B1(_1292_),
    .B2(_1285_),
    .A2(_1289_),
    .A1(_1284_));
 sg13g2_nor2b_1 _3625_ (.A(_1287_),
    .B_N(_1293_),
    .Y(_1294_));
 sg13g2_nand2_1 _3626_ (.Y(_1295_),
    .A(_1238_),
    .B(_1245_));
 sg13g2_nor4_1 _3627_ (.A(_1239_),
    .B(_1244_),
    .C(_1294_),
    .D(_1295_),
    .Y(_1296_));
 sg13g2_nor2_1 _3628_ (.A(net750),
    .B(_0662_),
    .Y(_1297_));
 sg13g2_a21oi_1 _3629_ (.A1(_1243_),
    .A2(_1296_),
    .Y(_1298_),
    .B1(_0662_));
 sg13g2_a21o_1 _3630_ (.A2(_1296_),
    .A1(_1243_),
    .B1(_0662_),
    .X(_1299_));
 sg13g2_nand2_2 _3631_ (.Y(_1300_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .B(_0647_));
 sg13g2_o21ai_1 _3632_ (.B1(net614),
    .Y(_1301_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .A2(net552));
 sg13g2_nor2_1 _3633_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .B(net585),
    .Y(_1302_));
 sg13g2_nand2b_2 _3634_ (.Y(_1303_),
    .B(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ));
 sg13g2_nor2_1 _3635_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .B(net567),
    .Y(_1304_));
 sg13g2_nor2_1 _3636_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .B(net573),
    .Y(_1305_));
 sg13g2_nor4_1 _3637_ (.A(_1301_),
    .B(_1302_),
    .C(_1304_),
    .D(_1305_),
    .Y(_1306_));
 sg13g2_o21ai_1 _3638_ (.B1(net597),
    .Y(_1307_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .A2(net559));
 sg13g2_nor2_1 _3639_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .B(net581),
    .Y(_1308_));
 sg13g2_nor2_1 _3640_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .B(net569),
    .Y(_1309_));
 sg13g2_nor2_1 _3641_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .B(net591),
    .Y(_1310_));
 sg13g2_nor4_1 _3642_ (.A(_1307_),
    .B(_1308_),
    .C(_1309_),
    .D(_1310_),
    .Y(_1311_));
 sg13g2_nor3_1 _3643_ (.A(net625),
    .B(_1306_),
    .C(_1311_),
    .Y(_1312_));
 sg13g2_o21ai_1 _3644_ (.B1(net597),
    .Y(_1313_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .A2(net591));
 sg13g2_nor2_1 _3645_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .B(net558),
    .Y(_1314_));
 sg13g2_nor2_1 _3646_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .B(net569),
    .Y(_1315_));
 sg13g2_nor2_1 _3647_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .B(net580),
    .Y(_1316_));
 sg13g2_nor4_1 _3648_ (.A(_1313_),
    .B(_1314_),
    .C(_1315_),
    .D(_1316_),
    .Y(_1317_));
 sg13g2_o21ai_1 _3649_ (.B1(net617),
    .Y(_1318_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .A2(net590));
 sg13g2_nor2_1 _3650_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .B(net568),
    .Y(_1319_));
 sg13g2_nor2_1 _3651_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .B(net558),
    .Y(_1320_));
 sg13g2_nor2_1 _3652_ (.A(_1319_),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_o21ai_1 _3653_ (.B1(_1321_),
    .Y(_1322_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .A2(net580));
 sg13g2_o21ai_1 _3654_ (.B1(net625),
    .Y(_1323_),
    .A1(_1318_),
    .A2(_1322_));
 sg13g2_o21ai_1 _3655_ (.B1(net613),
    .Y(_1324_),
    .A1(_1317_),
    .A2(_1323_));
 sg13g2_o21ai_1 _3656_ (.B1(net598),
    .Y(_1325_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .A2(net551));
 sg13g2_nor2_1 _3657_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .B(net562),
    .Y(_1326_));
 sg13g2_nor2_1 _3658_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .B(net574),
    .Y(_1327_));
 sg13g2_nor2_1 _3659_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .B(net585),
    .Y(_1328_));
 sg13g2_nor4_1 _3660_ (.A(_1325_),
    .B(_1326_),
    .C(_1327_),
    .D(_1328_),
    .Y(_1329_));
 sg13g2_o21ai_1 _3661_ (.B1(net614),
    .Y(_1330_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .A2(net561));
 sg13g2_nor2_1 _3662_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .B(net585),
    .Y(_1331_));
 sg13g2_nor2_1 _3663_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .B(net550),
    .Y(_1332_));
 sg13g2_nor2_1 _3664_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .B(net573),
    .Y(_1333_));
 sg13g2_nor4_1 _3665_ (.A(_1330_),
    .B(_1331_),
    .C(_1332_),
    .D(_1333_),
    .Y(_1334_));
 sg13g2_nor3_1 _3666_ (.A(_0646_),
    .B(_1329_),
    .C(_1334_),
    .Y(_1335_));
 sg13g2_o21ai_1 _3667_ (.B1(net614),
    .Y(_1336_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .A2(net584));
 sg13g2_nor2_1 _3668_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .B(net551),
    .Y(_1337_));
 sg13g2_nor2_1 _3669_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .B(net561),
    .Y(_1338_));
 sg13g2_nor2_1 _3670_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .B(net574),
    .Y(_1339_));
 sg13g2_nor4_1 _3671_ (.A(_1336_),
    .B(_1337_),
    .C(_1338_),
    .D(_1339_),
    .Y(_1340_));
 sg13g2_o21ai_1 _3672_ (.B1(net598),
    .Y(_1341_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .A2(net562));
 sg13g2_nor2_1 _3673_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .B(net586),
    .Y(_1342_));
 sg13g2_nor2_1 _3674_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .B(net575),
    .Y(_1343_));
 sg13g2_nor2_1 _3675_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .B(net550),
    .Y(_1344_));
 sg13g2_nor4_1 _3676_ (.A(_1341_),
    .B(_1342_),
    .C(_1343_),
    .D(_1344_),
    .Y(_1345_));
 sg13g2_nor3_1 _3677_ (.A(net618),
    .B(_1340_),
    .C(_1345_),
    .Y(_1346_));
 sg13g2_nor3_1 _3678_ (.A(net612),
    .B(_1335_),
    .C(_1346_),
    .Y(_1347_));
 sg13g2_nor2_1 _3679_ (.A(net610),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_o21ai_1 _3680_ (.B1(_1348_),
    .Y(_1349_),
    .A1(_1312_),
    .A2(_1324_));
 sg13g2_o21ai_1 _3681_ (.B1(net615),
    .Y(_1350_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .A2(net563));
 sg13g2_nor2_1 _3682_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .B(net586),
    .Y(_1351_));
 sg13g2_nor2_1 _3683_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .B(net575),
    .Y(_1352_));
 sg13g2_nor2_1 _3684_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .B(net553),
    .Y(_1353_));
 sg13g2_nor4_1 _3685_ (.A(_1350_),
    .B(_1351_),
    .C(_1352_),
    .D(_1353_),
    .Y(_1354_));
 sg13g2_o21ai_1 _3686_ (.B1(net597),
    .Y(_1355_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .A2(net580));
 sg13g2_nor2_1 _3687_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .B(net568),
    .Y(_1356_));
 sg13g2_nor2_1 _3688_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .B(net590),
    .Y(_1357_));
 sg13g2_nor2_1 _3689_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .B(net558),
    .Y(_1358_));
 sg13g2_nor4_1 _3690_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .D(_1358_),
    .Y(_1359_));
 sg13g2_nor3_1 _3691_ (.A(net625),
    .B(_1354_),
    .C(_1359_),
    .Y(_1360_));
 sg13g2_o21ai_1 _3692_ (.B1(net598),
    .Y(_1361_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .A2(net586));
 sg13g2_nor2_1 _3693_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .B(net564),
    .Y(_1362_));
 sg13g2_nor2_1 _3694_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .B(net554),
    .Y(_1363_));
 sg13g2_nor2_1 _3695_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .B(net576),
    .Y(_1364_));
 sg13g2_nor4_1 _3696_ (.A(_1361_),
    .B(_1362_),
    .C(_1363_),
    .D(_1364_),
    .Y(_1365_));
 sg13g2_o21ai_1 _3697_ (.B1(net615),
    .Y(_1366_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .A2(net564));
 sg13g2_nor2_1 _3698_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .B(net553),
    .Y(_1367_));
 sg13g2_a21oi_1 _3699_ (.A1(_0634_),
    .A2(net593),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_o21ai_1 _3700_ (.B1(_1368_),
    .Y(_1369_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .A2(net575));
 sg13g2_o21ai_1 _3701_ (.B1(net622),
    .Y(_1370_),
    .A1(_1366_),
    .A2(_1369_));
 sg13g2_o21ai_1 _3702_ (.B1(net612),
    .Y(_1371_),
    .A1(_1365_),
    .A2(_1370_));
 sg13g2_o21ai_1 _3703_ (.B1(net596),
    .Y(_1372_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .A2(net578));
 sg13g2_nor2_1 _3704_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .B(net556),
    .Y(_1373_));
 sg13g2_nor2_1 _3705_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .B(net588),
    .Y(_1374_));
 sg13g2_nor2_1 _3706_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .B(net566),
    .Y(_1375_));
 sg13g2_nor4_1 _3707_ (.A(_1372_),
    .B(_1373_),
    .C(_1374_),
    .D(_1375_),
    .Y(_1376_));
 sg13g2_o21ai_1 _3708_ (.B1(net616),
    .Y(_1377_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .A2(net588));
 sg13g2_nor2_1 _3709_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .B(net556),
    .Y(_1378_));
 sg13g2_nor2_1 _3710_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .B(net567),
    .Y(_1379_));
 sg13g2_nor2_1 _3711_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .B(net578),
    .Y(_1380_));
 sg13g2_nor4_1 _3712_ (.A(_1377_),
    .B(_1378_),
    .C(_1379_),
    .D(_1380_),
    .Y(_1381_));
 sg13g2_nor3_1 _3713_ (.A(_0646_),
    .B(_1376_),
    .C(_1381_),
    .Y(_1382_));
 sg13g2_o21ai_1 _3714_ (.B1(net616),
    .Y(_1383_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .A2(net579));
 sg13g2_nor2_1 _3715_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .B(net589),
    .Y(_1384_));
 sg13g2_nor2_1 _3716_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .B(net566),
    .Y(_1385_));
 sg13g2_nor2_1 _3717_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .B(net557),
    .Y(_1386_));
 sg13g2_nor4_1 _3718_ (.A(_1383_),
    .B(_1384_),
    .C(_1385_),
    .D(_1386_),
    .Y(_1387_));
 sg13g2_o21ai_1 _3719_ (.B1(net596),
    .Y(_1388_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .A2(net556));
 sg13g2_nor2_1 _3720_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .B(net567),
    .Y(_1389_));
 sg13g2_nor2_1 _3721_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .B(net573),
    .Y(_1390_));
 sg13g2_nor2_1 _3722_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .B(net588),
    .Y(_1391_));
 sg13g2_nor4_1 _3723_ (.A(_1388_),
    .B(_1389_),
    .C(_1390_),
    .D(_1391_),
    .Y(_1392_));
 sg13g2_nor3_1 _3724_ (.A(net623),
    .B(_1387_),
    .C(_1392_),
    .Y(_1393_));
 sg13g2_nor3_1 _3725_ (.A(net611),
    .B(_1382_),
    .C(_1393_),
    .Y(_1394_));
 sg13g2_nor2b_1 _3726_ (.A(_1394_),
    .B_N(net610),
    .Y(_1395_));
 sg13g2_o21ai_1 _3727_ (.B1(_1395_),
    .Y(_1396_),
    .A1(_1360_),
    .A2(_1371_));
 sg13g2_and2_1 _3728_ (.A(net2),
    .B(_1396_),
    .X(_1397_));
 sg13g2_a22oi_1 _3729_ (.Y(_1398_),
    .B1(_1349_),
    .B2(_1397_),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[2] ),
    .A1(_0661_));
 sg13g2_inv_1 _3730_ (.Y(_1399_),
    .A(_1398_));
 sg13g2_nor2_1 _3731_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .B(net591),
    .Y(_1400_));
 sg13g2_nor2_1 _3732_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .B(net580),
    .Y(_1401_));
 sg13g2_nor2_1 _3733_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .B(net559),
    .Y(_1402_));
 sg13g2_o21ai_1 _3734_ (.B1(net625),
    .Y(_1403_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .A2(net569));
 sg13g2_nor4_1 _3735_ (.A(_1400_),
    .B(_1401_),
    .C(_1402_),
    .D(_1403_),
    .Y(_1404_));
 sg13g2_nor2_1 _3736_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .B(net559),
    .Y(_1405_));
 sg13g2_nor2_1 _3737_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .B(net569),
    .Y(_1406_));
 sg13g2_nand2b_1 _3738_ (.Y(_1407_),
    .B(net594),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ));
 sg13g2_o21ai_1 _3739_ (.B1(_1407_),
    .Y(_1408_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .A2(net581));
 sg13g2_nor4_1 _3740_ (.A(net626),
    .B(_1405_),
    .C(_1406_),
    .D(_1408_),
    .Y(_1409_));
 sg13g2_nor3_1 _3741_ (.A(net617),
    .B(_1404_),
    .C(_1409_),
    .Y(_1410_));
 sg13g2_o21ai_1 _3742_ (.B1(net622),
    .Y(_1411_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .A2(net555));
 sg13g2_nor2_1 _3743_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .B(net580),
    .Y(_1412_));
 sg13g2_nor2_1 _3744_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .B(net568),
    .Y(_1413_));
 sg13g2_nor2_1 _3745_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .B(net590),
    .Y(_1414_));
 sg13g2_nor4_1 _3746_ (.A(_1411_),
    .B(_1412_),
    .C(_1413_),
    .D(_1414_),
    .Y(_1415_));
 sg13g2_nor2_1 _3747_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .B(net565),
    .Y(_1416_));
 sg13g2_nor2_1 _3748_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .B(net587),
    .Y(_1417_));
 sg13g2_nand2b_1 _3749_ (.Y(_1418_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ));
 sg13g2_o21ai_1 _3750_ (.B1(_1418_),
    .Y(_1419_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .A2(net555));
 sg13g2_nor4_1 _3751_ (.A(net622),
    .B(_1416_),
    .C(_1417_),
    .D(_1419_),
    .Y(_1420_));
 sg13g2_nor3_1 _3752_ (.A(net596),
    .B(_1415_),
    .C(_1420_),
    .Y(_1421_));
 sg13g2_nand2b_1 _3753_ (.Y(_1422_),
    .B(net613),
    .A_N(_1421_));
 sg13g2_nor2_1 _3754_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .B(net561),
    .Y(_1423_));
 sg13g2_nor2_1 _3755_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .B(net584),
    .Y(_1424_));
 sg13g2_nand2b_1 _3756_ (.Y(_1425_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ));
 sg13g2_o21ai_1 _3757_ (.B1(_1425_),
    .Y(_1426_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .A2(net550));
 sg13g2_nor4_1 _3758_ (.A(net618),
    .B(_1423_),
    .C(_1424_),
    .D(_1426_),
    .Y(_1427_));
 sg13g2_o21ai_1 _3759_ (.B1(net618),
    .Y(_1428_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .A2(net550));
 sg13g2_nor2_1 _3760_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .B(net584),
    .Y(_1429_));
 sg13g2_nor2_1 _3761_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .B(net561),
    .Y(_1430_));
 sg13g2_nor2_1 _3762_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .B(net574),
    .Y(_1431_));
 sg13g2_nor4_1 _3763_ (.A(_1428_),
    .B(_1429_),
    .C(_1430_),
    .D(_1431_),
    .Y(_1432_));
 sg13g2_nor3_1 _3764_ (.A(net598),
    .B(_1427_),
    .C(_1432_),
    .Y(_1433_));
 sg13g2_o21ai_1 _3765_ (.B1(net618),
    .Y(_1434_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .A2(net562));
 sg13g2_nor2_1 _3766_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .B(net584),
    .Y(_1435_));
 sg13g2_nor2_1 _3767_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .B(net551),
    .Y(_1436_));
 sg13g2_nor2_1 _3768_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .B(net574),
    .Y(_1437_));
 sg13g2_nor4_1 _3769_ (.A(_1434_),
    .B(_1435_),
    .C(_1436_),
    .D(_1437_),
    .Y(_1438_));
 sg13g2_nor2_1 _3770_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .B(net575),
    .Y(_1439_));
 sg13g2_nor2_1 _3771_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .B(net563),
    .Y(_1440_));
 sg13g2_nand2b_1 _3772_ (.Y(_1441_),
    .B(net593),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ));
 sg13g2_o21ai_1 _3773_ (.B1(_1441_),
    .Y(_1442_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .A2(net553));
 sg13g2_nor4_1 _3774_ (.A(net621),
    .B(_1439_),
    .C(_1440_),
    .D(_1442_),
    .Y(_1443_));
 sg13g2_nor3_1 _3775_ (.A(net614),
    .B(_1438_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_nor3_1 _3776_ (.A(net612),
    .B(_1433_),
    .C(_1444_),
    .Y(_1445_));
 sg13g2_nor2_1 _3777_ (.A(net610),
    .B(_1445_),
    .Y(_1446_));
 sg13g2_o21ai_1 _3778_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_1410_),
    .A2(_1422_));
 sg13g2_o21ai_1 _3779_ (.B1(net622),
    .Y(_1448_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .A2(net587));
 sg13g2_nor2_1 _3780_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .B(net576),
    .Y(_1449_));
 sg13g2_nor2_1 _3781_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .B(net564),
    .Y(_1450_));
 sg13g2_nor2_1 _3782_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .B(net554),
    .Y(_1451_));
 sg13g2_nor4_1 _3783_ (.A(_1448_),
    .B(_1449_),
    .C(_1450_),
    .D(_1451_),
    .Y(_1452_));
 sg13g2_nor2_1 _3784_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .B(net568),
    .Y(_1453_));
 sg13g2_nor2_1 _3785_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .B(net590),
    .Y(_1454_));
 sg13g2_nand2b_1 _3786_ (.Y(_1455_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ));
 sg13g2_o21ai_1 _3787_ (.B1(_1455_),
    .Y(_1456_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .A2(net558));
 sg13g2_nor4_1 _3788_ (.A(net625),
    .B(_1453_),
    .C(_1454_),
    .D(_1456_),
    .Y(_1457_));
 sg13g2_nor3_1 _3789_ (.A(net617),
    .B(_1452_),
    .C(_1457_),
    .Y(_1458_));
 sg13g2_nor2_1 _3790_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .B(net554),
    .Y(_1459_));
 sg13g2_nor2_1 _3791_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .B(net575),
    .Y(_1460_));
 sg13g2_or2_1 _3792_ (.X(_1461_),
    .B(net563),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ));
 sg13g2_o21ai_1 _3793_ (.B1(_1461_),
    .Y(_1462_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .A2(net586));
 sg13g2_nor4_1 _3794_ (.A(net621),
    .B(_1459_),
    .C(_1460_),
    .D(_1462_),
    .Y(_1463_));
 sg13g2_o21ai_1 _3795_ (.B1(net621),
    .Y(_1464_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .A2(net563));
 sg13g2_a22oi_1 _3796_ (.Y(_1465_),
    .B1(_0701_),
    .B2(_0650_),
    .A2(net593),
    .A1(_0635_));
 sg13g2_o21ai_1 _3797_ (.B1(_1465_),
    .Y(_1466_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .A2(net553));
 sg13g2_o21ai_1 _3798_ (.B1(net615),
    .Y(_1467_),
    .A1(_1464_),
    .A2(_1466_));
 sg13g2_o21ai_1 _3799_ (.B1(net612),
    .Y(_1468_),
    .A1(_1463_),
    .A2(_1467_));
 sg13g2_nor2_1 _3800_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .B(net557),
    .Y(_1469_));
 sg13g2_nor2_1 _3801_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .B(net579),
    .Y(_1470_));
 sg13g2_or2_1 _3802_ (.X(_1471_),
    .B(net566),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ));
 sg13g2_o21ai_1 _3803_ (.B1(_1471_),
    .Y(_1472_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .A2(net589));
 sg13g2_nor4_1 _3804_ (.A(net623),
    .B(_1469_),
    .C(_1470_),
    .D(_1472_),
    .Y(_1473_));
 sg13g2_o21ai_1 _3805_ (.B1(net624),
    .Y(_1474_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .A2(net567));
 sg13g2_nor2_1 _3806_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .B(net588),
    .Y(_1475_));
 sg13g2_nor2_1 _3807_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .B(net556),
    .Y(_1476_));
 sg13g2_nor2_1 _3808_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .B(net578),
    .Y(_1477_));
 sg13g2_nor4_1 _3809_ (.A(_1474_),
    .B(_1475_),
    .C(_1476_),
    .D(_1477_),
    .Y(_1478_));
 sg13g2_nor3_1 _3810_ (.A(net596),
    .B(_1473_),
    .C(_1478_),
    .Y(_1479_));
 sg13g2_nor2_1 _3811_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .B(net557),
    .Y(_1480_));
 sg13g2_nor2_1 _3812_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .B(net566),
    .Y(_1481_));
 sg13g2_nor2_1 _3813_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .B(net589),
    .Y(_1482_));
 sg13g2_o21ai_1 _3814_ (.B1(net624),
    .Y(_1483_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .A2(net578));
 sg13g2_nor4_1 _3815_ (.A(_1480_),
    .B(_1481_),
    .C(_1482_),
    .D(_1483_),
    .Y(_1484_));
 sg13g2_nor2_1 _3816_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .B(net567),
    .Y(_1485_));
 sg13g2_nand2b_1 _3817_ (.Y(_1486_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ));
 sg13g2_nor2_1 _3818_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .B(net588),
    .Y(_1487_));
 sg13g2_o21ai_1 _3819_ (.B1(_1486_),
    .Y(_1488_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .A2(net556));
 sg13g2_nor4_1 _3820_ (.A(net623),
    .B(_1485_),
    .C(_1487_),
    .D(_1488_),
    .Y(_1489_));
 sg13g2_nor3_1 _3821_ (.A(net616),
    .B(_1484_),
    .C(_1489_),
    .Y(_1490_));
 sg13g2_nor3_1 _3822_ (.A(net611),
    .B(_1479_),
    .C(_1490_),
    .Y(_1491_));
 sg13g2_nor2b_1 _3823_ (.A(_1491_),
    .B_N(net610),
    .Y(_1492_));
 sg13g2_o21ai_1 _3824_ (.B1(_1492_),
    .Y(_1493_),
    .A1(_1458_),
    .A2(_1468_));
 sg13g2_nand3_1 _3825_ (.B(_1447_),
    .C(_1493_),
    .A(net2),
    .Y(_1494_));
 sg13g2_o21ai_1 _3826_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_0660_),
    .A2(net2));
 sg13g2_nor2_1 _3827_ (.A(_1399_),
    .B(_1495_),
    .Y(_1496_));
 sg13g2_o21ai_1 _3828_ (.B1(net615),
    .Y(_1497_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .A2(net586));
 sg13g2_nor2_1 _3829_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .B(net553),
    .Y(_1498_));
 sg13g2_nor2_1 _3830_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .B(net575),
    .Y(_1499_));
 sg13g2_nor2_1 _3831_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .B(net564),
    .Y(_1500_));
 sg13g2_nor4_1 _3832_ (.A(_1497_),
    .B(_1498_),
    .C(_1499_),
    .D(_1500_),
    .Y(_1501_));
 sg13g2_o21ai_1 _3833_ (.B1(net598),
    .Y(_1502_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .A2(net576));
 sg13g2_nor2_1 _3834_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .B(net590),
    .Y(_1503_));
 sg13g2_nor2_1 _3835_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .B(net558),
    .Y(_1504_));
 sg13g2_nor2_1 _3836_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .B(net568),
    .Y(_1505_));
 sg13g2_nor4_1 _3837_ (.A(_1502_),
    .B(_1503_),
    .C(_1504_),
    .D(_1505_),
    .Y(_1506_));
 sg13g2_nor3_1 _3838_ (.A(net622),
    .B(_1501_),
    .C(_1506_),
    .Y(_1507_));
 sg13g2_o21ai_1 _3839_ (.B1(net598),
    .Y(_1508_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .A2(net587));
 sg13g2_nor2_1 _3840_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .B(net576),
    .Y(_1509_));
 sg13g2_nor2_1 _3841_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .B(net554),
    .Y(_1510_));
 sg13g2_nor2_1 _3842_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .B(net565),
    .Y(_1511_));
 sg13g2_nor4_1 _3843_ (.A(_1508_),
    .B(_1509_),
    .C(_1510_),
    .D(_1511_),
    .Y(_1512_));
 sg13g2_o21ai_1 _3844_ (.B1(net615),
    .Y(_1513_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .A2(net553));
 sg13g2_nor2_1 _3845_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .B(net563),
    .Y(_1514_));
 sg13g2_a21oi_1 _3846_ (.A1(_0649_),
    .A2(_0701_),
    .Y(_1515_),
    .B1(_1514_));
 sg13g2_o21ai_1 _3847_ (.B1(_1515_),
    .Y(_1516_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .A2(net586));
 sg13g2_o21ai_1 _3848_ (.B1(net621),
    .Y(_1517_),
    .A1(_1513_),
    .A2(_1516_));
 sg13g2_o21ai_1 _3849_ (.B1(net612),
    .Y(_1518_),
    .A1(_1512_),
    .A2(_1517_));
 sg13g2_or2_1 _3850_ (.X(_1519_),
    .B(_1518_),
    .A(_1507_));
 sg13g2_o21ai_1 _3851_ (.B1(net596),
    .Y(_1520_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .A2(net566));
 sg13g2_nor2_1 _3852_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .B(net578),
    .Y(_1521_));
 sg13g2_nor2_1 _3853_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .B(net557),
    .Y(_1522_));
 sg13g2_nor2_1 _3854_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .B(net588),
    .Y(_1523_));
 sg13g2_nor4_1 _3855_ (.A(_1520_),
    .B(_1521_),
    .C(_1522_),
    .D(_1523_),
    .Y(_1524_));
 sg13g2_o21ai_1 _3856_ (.B1(net616),
    .Y(_1525_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .A2(net570));
 sg13g2_a22oi_1 _3857_ (.Y(_1526_),
    .B1(net583),
    .B2(_0633_),
    .A2(net594),
    .A1(_0632_));
 sg13g2_o21ai_1 _3858_ (.B1(_1526_),
    .Y(_1527_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .A2(net556));
 sg13g2_o21ai_1 _3859_ (.B1(net624),
    .Y(_1528_),
    .A1(_1525_),
    .A2(_1527_));
 sg13g2_nor2_1 _3860_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .B(net589),
    .Y(_1529_));
 sg13g2_nor2_1 _3861_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .B(net579),
    .Y(_1530_));
 sg13g2_o21ai_1 _3862_ (.B1(net616),
    .Y(_1531_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .A2(net557));
 sg13g2_nor3_1 _3863_ (.A(_1529_),
    .B(_1530_),
    .C(_1531_),
    .Y(_1532_));
 sg13g2_o21ai_1 _3864_ (.B1(_1532_),
    .Y(_1533_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .A2(net566));
 sg13g2_nor2_1 _3865_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .B(net567),
    .Y(_1534_));
 sg13g2_nor2_1 _3866_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .B(net573),
    .Y(_1535_));
 sg13g2_nor2_1 _3867_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .B(net585),
    .Y(_1536_));
 sg13g2_o21ai_1 _3868_ (.B1(net596),
    .Y(_1537_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .A2(net556));
 sg13g2_nor4_1 _3869_ (.A(_1534_),
    .B(_1535_),
    .C(_1536_),
    .D(_1537_),
    .Y(_1538_));
 sg13g2_nor2_1 _3870_ (.A(net624),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_a21oi_1 _3871_ (.A1(_1533_),
    .A2(_1539_),
    .Y(_1540_),
    .B1(net611));
 sg13g2_o21ai_1 _3872_ (.B1(_1540_),
    .Y(_1541_),
    .A1(_1524_),
    .A2(_1528_));
 sg13g2_nand3_1 _3873_ (.B(_1519_),
    .C(_1541_),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .Y(_1542_));
 sg13g2_o21ai_1 _3874_ (.B1(net620),
    .Y(_1543_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .A2(net584));
 sg13g2_nor2_1 _3875_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .B(net574),
    .Y(_1544_));
 sg13g2_nor2_1 _3876_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .B(net551),
    .Y(_1545_));
 sg13g2_nor2_1 _3877_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .B(net562),
    .Y(_1546_));
 sg13g2_nor4_1 _3878_ (.A(_1543_),
    .B(_1544_),
    .C(_1545_),
    .D(_1546_),
    .Y(_1547_));
 sg13g2_nor2_1 _3879_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .B(net563),
    .Y(_1548_));
 sg13g2_nor2_1 _3880_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .B(net586),
    .Y(_1549_));
 sg13g2_nand2b_1 _3881_ (.Y(_1550_),
    .B(_0701_),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ));
 sg13g2_o21ai_1 _3882_ (.B1(_1550_),
    .Y(_1551_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .A2(net553));
 sg13g2_nor4_1 _3883_ (.A(net621),
    .B(_1548_),
    .C(_1549_),
    .D(_1551_),
    .Y(_1552_));
 sg13g2_nor3_1 _3884_ (.A(net614),
    .B(_1547_),
    .C(_1552_),
    .Y(_1553_));
 sg13g2_o21ai_1 _3885_ (.B1(net618),
    .Y(_1554_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .A2(net561));
 sg13g2_nor2_1 _3886_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .B(net584),
    .Y(_1555_));
 sg13g2_nor2_1 _3887_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .B(net573),
    .Y(_1556_));
 sg13g2_nor2_1 _3888_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .B(net550),
    .Y(_1557_));
 sg13g2_nor4_1 _3889_ (.A(_1554_),
    .B(_1555_),
    .C(_1556_),
    .D(_1557_),
    .Y(_1558_));
 sg13g2_nor2_1 _3890_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .B(net574),
    .Y(_1559_));
 sg13g2_nor2_1 _3891_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .B(net550),
    .Y(_1560_));
 sg13g2_nand2b_1 _3892_ (.Y(_1561_),
    .B(net593),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ));
 sg13g2_o21ai_1 _3893_ (.B1(_1561_),
    .Y(_1562_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .A2(net561));
 sg13g2_nor4_1 _3894_ (.A(net618),
    .B(_1559_),
    .C(_1560_),
    .D(_1562_),
    .Y(_1563_));
 sg13g2_nor3_1 _3895_ (.A(net598),
    .B(_1558_),
    .C(_1563_),
    .Y(_1564_));
 sg13g2_nor3_1 _3896_ (.A(net612),
    .B(_1553_),
    .C(_1564_),
    .Y(_1565_));
 sg13g2_nor2_1 _3897_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .B(net591),
    .Y(_1566_));
 sg13g2_nor2_1 _3898_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .B(net569),
    .Y(_1567_));
 sg13g2_nor2_1 _3899_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .B(net581),
    .Y(_1568_));
 sg13g2_o21ai_1 _3900_ (.B1(net626),
    .Y(_1569_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .A2(net559));
 sg13g2_nor4_1 _3901_ (.A(_1566_),
    .B(_1567_),
    .C(_1568_),
    .D(_1569_),
    .Y(_1570_));
 sg13g2_nor2_1 _3902_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .B(net581),
    .Y(_1571_));
 sg13g2_nor2_1 _3903_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .B(net559),
    .Y(_1572_));
 sg13g2_nand2b_1 _3904_ (.Y(_1573_),
    .B(net594),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ));
 sg13g2_o21ai_1 _3905_ (.B1(_1573_),
    .Y(_1574_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .A2(net569));
 sg13g2_nor4_1 _3906_ (.A(net626),
    .B(_1571_),
    .C(_1572_),
    .D(_1574_),
    .Y(_1575_));
 sg13g2_nor3_1 _3907_ (.A(net616),
    .B(_1570_),
    .C(_1575_),
    .Y(_1576_));
 sg13g2_o21ai_1 _3908_ (.B1(net625),
    .Y(_1577_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .A2(net590));
 sg13g2_nor2_1 _3909_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .B(net580),
    .Y(_1578_));
 sg13g2_nor2_1 _3910_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .B(net558),
    .Y(_1579_));
 sg13g2_nor2_1 _3911_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .B(net568),
    .Y(_1580_));
 sg13g2_nor4_1 _3912_ (.A(_1577_),
    .B(_1578_),
    .C(_1579_),
    .D(_1580_),
    .Y(_1581_));
 sg13g2_nor2_1 _3913_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .B(net552),
    .Y(_1582_));
 sg13g2_nand2b_1 _3914_ (.Y(_1583_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ));
 sg13g2_o21ai_1 _3915_ (.B1(_1583_),
    .Y(_1584_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .A2(net585));
 sg13g2_nor2_1 _3916_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .B(net565),
    .Y(_1585_));
 sg13g2_nor4_1 _3917_ (.A(net619),
    .B(_1582_),
    .C(_1584_),
    .D(_1585_),
    .Y(_1586_));
 sg13g2_nor3_1 _3918_ (.A(net597),
    .B(_1581_),
    .C(_1586_),
    .Y(_1587_));
 sg13g2_nor3_1 _3919_ (.A(_0644_),
    .B(_1576_),
    .C(_1587_),
    .Y(_1588_));
 sg13g2_nor3_1 _3920_ (.A(net610),
    .B(_1565_),
    .C(_1588_),
    .Y(_1589_));
 sg13g2_nor2_1 _3921_ (.A(_0661_),
    .B(_1589_),
    .Y(_1590_));
 sg13g2_a22oi_1 _3922_ (.Y(_1591_),
    .B1(_1542_),
    .B2(_1590_),
    .A2(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .A1(_0661_));
 sg13g2_nor2_1 _3923_ (.A(net749),
    .B(net1),
    .Y(_1592_));
 sg13g2_nor2_1 _3924_ (.A(net1),
    .B(_1591_),
    .Y(_1593_));
 sg13g2_nand2_1 _3925_ (.Y(_1594_),
    .A(net797),
    .B(_1593_));
 sg13g2_nor2_1 _3926_ (.A(_1496_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_a21oi_1 _3927_ (.A1(net797),
    .A2(_1298_),
    .Y(_1596_),
    .B1(_1595_));
 sg13g2_inv_1 _3928_ (.Y(_0372_),
    .A(_1596_));
 sg13g2_o21ai_1 _3929_ (.B1(net626),
    .Y(_1597_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .A2(net581));
 sg13g2_nor2_1 _3930_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .B(net591),
    .Y(_1598_));
 sg13g2_nor2_1 _3931_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .B(net559),
    .Y(_1599_));
 sg13g2_nor2_1 _3932_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .B(net569),
    .Y(_1600_));
 sg13g2_nor4_1 _3933_ (.A(_1597_),
    .B(_1598_),
    .C(_1599_),
    .D(_1600_),
    .Y(_1601_));
 sg13g2_nor2_1 _3934_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .B(net581),
    .Y(_1602_));
 sg13g2_nor2_1 _3935_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .B(net569),
    .Y(_1603_));
 sg13g2_nand2b_1 _3936_ (.Y(_1604_),
    .B(net594),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ));
 sg13g2_o21ai_1 _3937_ (.B1(_1604_),
    .Y(_1605_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .A2(net559));
 sg13g2_nor4_1 _3938_ (.A(net626),
    .B(_1602_),
    .C(_1603_),
    .D(_1605_),
    .Y(_1606_));
 sg13g2_nor3_1 _3939_ (.A(net617),
    .B(_1601_),
    .C(_1606_),
    .Y(_1607_));
 sg13g2_o21ai_1 _3940_ (.B1(net625),
    .Y(_1608_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .A2(net590));
 sg13g2_nor2_1 _3941_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ),
    .B(net580),
    .Y(_1609_));
 sg13g2_nor2_1 _3942_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .B(net568),
    .Y(_1610_));
 sg13g2_nor2_1 _3943_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ),
    .B(net558),
    .Y(_1611_));
 sg13g2_nor4_1 _3944_ (.A(_1608_),
    .B(_1609_),
    .C(_1610_),
    .D(_1611_),
    .Y(_1612_));
 sg13g2_nor2_1 _3945_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .B(net564),
    .Y(_1613_));
 sg13g2_nand2b_1 _3946_ (.Y(_1614_),
    .B(net593),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ));
 sg13g2_o21ai_1 _3947_ (.B1(_1614_),
    .Y(_1615_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .A2(net577));
 sg13g2_nor2_1 _3948_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ),
    .B(net555),
    .Y(_1616_));
 sg13g2_nor4_1 _3949_ (.A(net622),
    .B(_1613_),
    .C(_1615_),
    .D(_1616_),
    .Y(_1617_));
 sg13g2_nor3_1 _3950_ (.A(net597),
    .B(_1612_),
    .C(_1617_),
    .Y(_1618_));
 sg13g2_nand2b_1 _3951_ (.Y(_1619_),
    .B(net613),
    .A_N(_1618_));
 sg13g2_nor2_1 _3952_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .B(net574),
    .Y(_1620_));
 sg13g2_nor2_1 _3953_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .B(net550),
    .Y(_1621_));
 sg13g2_nand2b_1 _3954_ (.Y(_1622_),
    .B(net593),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ));
 sg13g2_o21ai_1 _3955_ (.B1(_1622_),
    .Y(_1623_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .A2(net561));
 sg13g2_nor4_1 _3956_ (.A(net618),
    .B(_1620_),
    .C(_1621_),
    .D(_1623_),
    .Y(_1624_));
 sg13g2_o21ai_1 _3957_ (.B1(net618),
    .Y(_1625_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .A2(net550));
 sg13g2_nor2_1 _3958_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .B(net561),
    .Y(_1626_));
 sg13g2_nor2_1 _3959_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .B(net573),
    .Y(_1627_));
 sg13g2_nor2_1 _3960_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .B(net584),
    .Y(_1628_));
 sg13g2_nor4_1 _3961_ (.A(_1625_),
    .B(_1626_),
    .C(_1627_),
    .D(_1628_),
    .Y(_1629_));
 sg13g2_nor3_1 _3962_ (.A(net598),
    .B(_1624_),
    .C(_1629_),
    .Y(_1630_));
 sg13g2_o21ai_1 _3963_ (.B1(net620),
    .Y(_1631_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .A2(net574));
 sg13g2_nor2_1 _3964_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .B(net562),
    .Y(_1632_));
 sg13g2_nor2_1 _3965_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .B(net551),
    .Y(_1633_));
 sg13g2_nor2_1 _3966_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .B(net584),
    .Y(_1634_));
 sg13g2_nor4_1 _3967_ (.A(_1631_),
    .B(_1632_),
    .C(_1633_),
    .D(_1634_),
    .Y(_1635_));
 sg13g2_nor2_1 _3968_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .B(net563),
    .Y(_1636_));
 sg13g2_nor2_1 _3969_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .B(net575),
    .Y(_1637_));
 sg13g2_nand2b_1 _3970_ (.Y(_1638_),
    .B(net594),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ));
 sg13g2_o21ai_1 _3971_ (.B1(_1638_),
    .Y(_1639_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .A2(net553));
 sg13g2_nor4_1 _3972_ (.A(net621),
    .B(_1636_),
    .C(_1637_),
    .D(_1639_),
    .Y(_1640_));
 sg13g2_nor3_1 _3973_ (.A(net614),
    .B(_1635_),
    .C(_1640_),
    .Y(_1641_));
 sg13g2_nor3_2 _3974_ (.A(net612),
    .B(_1630_),
    .C(_1641_),
    .Y(_1642_));
 sg13g2_nor2_1 _3975_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_o21ai_1 _3976_ (.B1(_1643_),
    .Y(_1644_),
    .A1(_1607_),
    .A2(_1619_));
 sg13g2_o21ai_1 _3977_ (.B1(net622),
    .Y(_1645_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ),
    .A2(net576));
 sg13g2_nor2_1 _3978_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .B(net554),
    .Y(_1646_));
 sg13g2_nor2_1 _3979_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ),
    .B(net586),
    .Y(_1647_));
 sg13g2_nor2_1 _3980_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .B(net564),
    .Y(_1648_));
 sg13g2_nor4_1 _3981_ (.A(_1645_),
    .B(_1646_),
    .C(_1647_),
    .D(_1648_),
    .Y(_1649_));
 sg13g2_nor2_1 _3982_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .B(net590),
    .Y(_1650_));
 sg13g2_nor2_1 _3983_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .B(net580),
    .Y(_1651_));
 sg13g2_or2_1 _3984_ (.X(_1652_),
    .B(net568),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ));
 sg13g2_o21ai_1 _3985_ (.B1(_1652_),
    .Y(_1653_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .A2(net558));
 sg13g2_nor4_1 _3986_ (.A(net625),
    .B(_1650_),
    .C(_1651_),
    .D(_1653_),
    .Y(_1654_));
 sg13g2_nor3_1 _3987_ (.A(net617),
    .B(_1649_),
    .C(_1654_),
    .Y(_1655_));
 sg13g2_nor2_1 _3988_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .B(net564),
    .Y(_1656_));
 sg13g2_nor2_1 _3989_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .B(net576),
    .Y(_1657_));
 sg13g2_nand2b_1 _3990_ (.Y(_1658_),
    .B(net594),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ));
 sg13g2_o21ai_1 _3991_ (.B1(_1658_),
    .Y(_1659_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .A2(net554));
 sg13g2_nor4_1 _3992_ (.A(net621),
    .B(_1656_),
    .C(_1657_),
    .D(_1659_),
    .Y(_1660_));
 sg13g2_o21ai_1 _3993_ (.B1(net621),
    .Y(_1661_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .A2(net575));
 sg13g2_nor2_1 _3994_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .B(net563),
    .Y(_1662_));
 sg13g2_a21oi_1 _3995_ (.A1(_0636_),
    .A2(net594),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_o21ai_1 _3996_ (.B1(_1663_),
    .Y(_1664_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .A2(net554));
 sg13g2_o21ai_1 _3997_ (.B1(net615),
    .Y(_1665_),
    .A1(_1661_),
    .A2(_1664_));
 sg13g2_o21ai_1 _3998_ (.B1(net612),
    .Y(_1666_),
    .A1(_1660_),
    .A2(_1665_));
 sg13g2_or2_1 _3999_ (.X(_1667_),
    .B(_1666_),
    .A(_1655_));
 sg13g2_nor2_1 _4000_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .B(net589),
    .Y(_1668_));
 sg13g2_nor2_1 _4001_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .B(net557),
    .Y(_1669_));
 sg13g2_or2_1 _4002_ (.X(_1670_),
    .B(net566),
    .A(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ));
 sg13g2_o21ai_1 _4003_ (.B1(_1670_),
    .Y(_1671_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .A2(net579));
 sg13g2_nor4_1 _4004_ (.A(net623),
    .B(_1668_),
    .C(_1669_),
    .D(_1671_),
    .Y(_1672_));
 sg13g2_o21ai_1 _4005_ (.B1(net624),
    .Y(_1673_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ),
    .A2(net570));
 sg13g2_nor2_1 _4006_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .B(net588),
    .Y(_1674_));
 sg13g2_nor2_1 _4007_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ),
    .B(net557),
    .Y(_1675_));
 sg13g2_nor2_1 _4008_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .B(net578),
    .Y(_1676_));
 sg13g2_nor4_1 _4009_ (.A(_1673_),
    .B(_1674_),
    .C(_1675_),
    .D(_1676_),
    .Y(_1677_));
 sg13g2_nor3_1 _4010_ (.A(net596),
    .B(_1672_),
    .C(_1677_),
    .Y(_1678_));
 sg13g2_nor2_1 _4011_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .B(net589),
    .Y(_1679_));
 sg13g2_nor2_1 _4012_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .B(net557),
    .Y(_1680_));
 sg13g2_nor2_1 _4013_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .B(net579),
    .Y(_1681_));
 sg13g2_o21ai_1 _4014_ (.B1(net623),
    .Y(_1682_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .A2(net566));
 sg13g2_nor4_1 _4015_ (.A(_1679_),
    .B(_1680_),
    .C(_1681_),
    .D(_1682_),
    .Y(_1683_));
 sg13g2_nor2_1 _4016_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .B(net567),
    .Y(_1684_));
 sg13g2_nor2_1 _4017_ (.A(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .B(net556),
    .Y(_1685_));
 sg13g2_nand2b_1 _4018_ (.Y(_1686_),
    .B(net583),
    .A_N(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ));
 sg13g2_o21ai_1 _4019_ (.B1(_1686_),
    .Y(_1687_),
    .A1(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .A2(net588));
 sg13g2_nor4_1 _4020_ (.A(net623),
    .B(_1684_),
    .C(_1685_),
    .D(_1687_),
    .Y(_1688_));
 sg13g2_nor3_1 _4021_ (.A(net616),
    .B(_1683_),
    .C(_1688_),
    .Y(_1689_));
 sg13g2_nor3_1 _4022_ (.A(net611),
    .B(_1678_),
    .C(_1689_),
    .Y(_1690_));
 sg13g2_nor2b_1 _4023_ (.A(_1690_),
    .B_N(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .Y(_1691_));
 sg13g2_a21oi_1 _4024_ (.A1(_1667_),
    .A2(_1691_),
    .Y(_1692_),
    .B1(_0661_));
 sg13g2_a22oi_1 _4025_ (.Y(_1693_),
    .B1(_1644_),
    .B2(_1692_),
    .A2(_0661_),
    .A1(\videogen.test_lut_thingy.gol_counter_reg[0] ));
 sg13g2_inv_1 _4026_ (.Y(_1694_),
    .A(_1693_));
 sg13g2_nand2_1 _4027_ (.Y(_1695_),
    .A(_1495_),
    .B(_1693_));
 sg13g2_inv_1 _4028_ (.Y(_1696_),
    .A(_1695_));
 sg13g2_a21oi_1 _4029_ (.A1(_1299_),
    .A2(_1696_),
    .Y(_0374_),
    .B1(_1596_));
 sg13g2_nor2b_1 _4030_ (.A(_1398_),
    .B_N(_1495_),
    .Y(_1697_));
 sg13g2_nor2_1 _4031_ (.A(_1398_),
    .B(_1695_),
    .Y(_1698_));
 sg13g2_a21oi_1 _4032_ (.A1(_1299_),
    .A2(_1698_),
    .Y(_0373_),
    .B1(_1596_));
 sg13g2_nand2b_1 _4033_ (.Y(_1699_),
    .B(_1693_),
    .A_N(_1495_));
 sg13g2_inv_1 _4034_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_a21oi_1 _4035_ (.A1(_1398_),
    .A2(_1700_),
    .Y(_1701_),
    .B1(_1594_));
 sg13g2_a21o_1 _4036_ (.A2(_1298_),
    .A1(net798),
    .B1(_1701_),
    .X(_0375_));
 sg13g2_o21ai_1 _4037_ (.B1(_0990_),
    .Y(_1702_),
    .A1(_0989_),
    .A2(_1059_));
 sg13g2_xnor2_1 _4038_ (.Y(_1703_),
    .A(_1060_),
    .B(_1702_));
 sg13g2_xnor2_1 _4039_ (.Y(_1704_),
    .A(_0995_),
    .B(_1195_));
 sg13g2_inv_1 _4040_ (.Y(_1705_),
    .A(_1704_));
 sg13g2_nand2_2 _4041_ (.Y(_1706_),
    .A(_0995_),
    .B(_1192_));
 sg13g2_xnor2_1 _4042_ (.Y(_1707_),
    .A(_1076_),
    .B(_1706_));
 sg13g2_nor2_1 _4043_ (.A(_1073_),
    .B(_1706_),
    .Y(_1708_));
 sg13g2_nor2_1 _4044_ (.A(_1093_),
    .B(_1706_),
    .Y(_1709_));
 sg13g2_and2_1 _4045_ (.A(_1100_),
    .B(_1709_),
    .X(_1710_));
 sg13g2_or3_1 _4046_ (.A(_1164_),
    .B(_1165_),
    .C(_1710_),
    .X(_1711_));
 sg13g2_o21ai_1 _4047_ (.B1(_1710_),
    .Y(_1712_),
    .A1(_1164_),
    .A2(_1165_));
 sg13g2_nand2_1 _4048_ (.Y(_1713_),
    .A(_1711_),
    .B(_1712_));
 sg13g2_and2_1 _4049_ (.A(_1145_),
    .B(_1709_),
    .X(_1714_));
 sg13g2_or3_1 _4050_ (.A(_1156_),
    .B(_1157_),
    .C(_1714_),
    .X(_1715_));
 sg13g2_o21ai_1 _4051_ (.B1(_1714_),
    .Y(_1716_),
    .A1(_1156_),
    .A2(_1157_));
 sg13g2_nand2_2 _4052_ (.Y(_1717_),
    .A(_1715_),
    .B(_1716_));
 sg13g2_xnor2_1 _4053_ (.Y(_1718_),
    .A(_1147_),
    .B(_1709_));
 sg13g2_a221oi_1 _4054_ (.B2(_1716_),
    .C1(_1718_),
    .B1(_1715_),
    .A1(_1711_),
    .Y(_1719_),
    .A2(_1712_));
 sg13g2_and2_1 _4055_ (.A(_1163_),
    .B(_1710_),
    .X(_1720_));
 sg13g2_a21oi_2 _4056_ (.B1(_1720_),
    .Y(_1721_),
    .A2(_1137_),
    .A1(_1135_));
 sg13g2_and3_2 _4057_ (.X(_1722_),
    .A(_1135_),
    .B(_1137_),
    .C(_1720_));
 sg13g2_nor2_2 _4058_ (.A(_1721_),
    .B(_1722_),
    .Y(_1723_));
 sg13g2_nor4_1 _4059_ (.A(_1718_),
    .B(_1719_),
    .C(_1721_),
    .D(_1722_),
    .Y(_1724_));
 sg13g2_or4_1 _4060_ (.A(_1718_),
    .B(_1719_),
    .C(_1721_),
    .D(_1722_),
    .X(_1725_));
 sg13g2_a21o_1 _4061_ (.A2(_1724_),
    .A1(_1717_),
    .B1(_1713_),
    .X(_1726_));
 sg13g2_o21ai_1 _4062_ (.B1(_1718_),
    .Y(_1727_),
    .A1(_1721_),
    .A2(_1722_));
 sg13g2_and2_1 _4063_ (.A(_1725_),
    .B(_1727_),
    .X(_1728_));
 sg13g2_xnor2_1 _4064_ (.Y(_1729_),
    .A(net544),
    .B(_1708_));
 sg13g2_and4_1 _4065_ (.A(_1717_),
    .B(_1725_),
    .C(_1727_),
    .D(_1729_),
    .X(_1730_));
 sg13g2_nand2_1 _4066_ (.Y(_1731_),
    .A(_1719_),
    .B(_1723_));
 sg13g2_o21ai_1 _4067_ (.B1(_1731_),
    .Y(_1732_),
    .A1(_1726_),
    .A2(_1730_));
 sg13g2_o21ai_1 _4068_ (.B1(_1726_),
    .Y(_1733_),
    .A1(_1730_),
    .A2(_1731_));
 sg13g2_o21ai_1 _4069_ (.B1(_1733_),
    .Y(_1734_),
    .A1(_1726_),
    .A2(_1730_));
 sg13g2_xnor2_1 _4070_ (.Y(_1735_),
    .A(_1717_),
    .B(_1724_));
 sg13g2_nand2_1 _4071_ (.Y(_1736_),
    .A(_1729_),
    .B(_1732_));
 sg13g2_nand3_1 _4072_ (.B(_1729_),
    .C(_1732_),
    .A(_1728_),
    .Y(_1737_));
 sg13g2_a22oi_1 _4073_ (.Y(_1738_),
    .B1(_1735_),
    .B2(_1737_),
    .A2(_1732_),
    .A1(_1730_));
 sg13g2_xor2_1 _4074_ (.B(_1732_),
    .A(_1729_),
    .X(_1739_));
 sg13g2_and3_1 _4075_ (.X(_1740_),
    .A(_1707_),
    .B(_1728_),
    .C(_1739_));
 sg13g2_nor2_1 _4076_ (.A(_1738_),
    .B(_1740_),
    .Y(_1741_));
 sg13g2_o21ai_1 _4077_ (.B1(_1734_),
    .Y(_1742_),
    .A1(_1738_),
    .A2(_1740_));
 sg13g2_nand2_1 _4078_ (.Y(_1743_),
    .A(_1707_),
    .B(_1742_));
 sg13g2_inv_1 _4079_ (.Y(_1744_),
    .A(_1743_));
 sg13g2_xnor2_1 _4080_ (.Y(_1745_),
    .A(_1707_),
    .B(_1742_));
 sg13g2_nand2_1 _4081_ (.Y(_1746_),
    .A(_1704_),
    .B(_1739_));
 sg13g2_or2_1 _4082_ (.X(_1747_),
    .B(_1746_),
    .A(_1745_));
 sg13g2_xor2_1 _4083_ (.B(_1736_),
    .A(_1728_),
    .X(_1748_));
 sg13g2_nand3_1 _4084_ (.B(_1739_),
    .C(_1742_),
    .A(_1707_),
    .Y(_1749_));
 sg13g2_xnor2_1 _4085_ (.Y(_1750_),
    .A(_1748_),
    .B(_1749_));
 sg13g2_o21ai_1 _4086_ (.B1(_1738_),
    .Y(_1751_),
    .A1(_1734_),
    .A2(_1740_));
 sg13g2_nor2b_1 _4087_ (.A(_1741_),
    .B_N(_1751_),
    .Y(_1752_));
 sg13g2_a21oi_1 _4088_ (.A1(_1747_),
    .A2(_1750_),
    .Y(_1753_),
    .B1(_1752_));
 sg13g2_xnor2_1 _4089_ (.Y(_1754_),
    .A(_1705_),
    .B(_1753_));
 sg13g2_nand2b_1 _4090_ (.Y(_1755_),
    .B(_1065_),
    .A_N(_0990_));
 sg13g2_nand2_1 _4091_ (.Y(_1756_),
    .A(_0990_),
    .B(_1066_));
 sg13g2_and2_1 _4092_ (.A(_1755_),
    .B(_1756_),
    .X(_1757_));
 sg13g2_nor3_1 _4093_ (.A(_1745_),
    .B(_1754_),
    .C(_1757_),
    .Y(_1758_));
 sg13g2_nor3_1 _4094_ (.A(_1705_),
    .B(_1745_),
    .C(_1753_),
    .Y(_1759_));
 sg13g2_or3_1 _4095_ (.A(_1739_),
    .B(_1744_),
    .C(_1759_),
    .X(_1760_));
 sg13g2_o21ai_1 _4096_ (.B1(_1739_),
    .Y(_1761_),
    .A1(_1744_),
    .A2(_1759_));
 sg13g2_and2_1 _4097_ (.A(_1760_),
    .B(_1761_),
    .X(_1762_));
 sg13g2_a21o_1 _4098_ (.A2(_1761_),
    .A1(_1760_),
    .B1(_1758_),
    .X(_1763_));
 sg13g2_a21oi_1 _4099_ (.A1(_1747_),
    .A2(_1752_),
    .Y(_1764_),
    .B1(_1750_));
 sg13g2_a21o_2 _4100_ (.A2(_1750_),
    .A1(_1747_),
    .B1(_1764_),
    .X(_1765_));
 sg13g2_o21ai_1 _4101_ (.B1(_1762_),
    .Y(_1766_),
    .A1(_1758_),
    .A2(_1765_));
 sg13g2_and2_1 _4102_ (.A(_1763_),
    .B(_1766_),
    .X(_1767_));
 sg13g2_a21oi_1 _4103_ (.A1(_1763_),
    .A2(_1765_),
    .Y(_1768_),
    .B1(_1757_));
 sg13g2_nand3_1 _4104_ (.B(_1762_),
    .C(_1765_),
    .A(_1757_),
    .Y(_1769_));
 sg13g2_nand2b_1 _4105_ (.Y(_1770_),
    .B(_1769_),
    .A_N(_1768_));
 sg13g2_nor2_1 _4106_ (.A(_1703_),
    .B(_1754_),
    .Y(_1771_));
 sg13g2_nand3b_1 _4107_ (.B(_1769_),
    .C(_1771_),
    .Y(_1772_),
    .A_N(_1768_));
 sg13g2_a221oi_1 _4108_ (.B2(_1765_),
    .C1(_1754_),
    .B1(_1763_),
    .A1(_1755_),
    .Y(_1773_),
    .A2(_1756_));
 sg13g2_o21ai_1 _4109_ (.B1(_1745_),
    .Y(_1774_),
    .A1(_1705_),
    .A2(_1753_));
 sg13g2_nor2b_1 _4110_ (.A(_1759_),
    .B_N(_1774_),
    .Y(_1775_));
 sg13g2_xnor2_1 _4111_ (.Y(_1776_),
    .A(_1773_),
    .B(_1775_));
 sg13g2_a21oi_2 _4112_ (.B1(_1767_),
    .Y(_1777_),
    .A2(_1776_),
    .A1(_1772_));
 sg13g2_xor2_1 _4113_ (.B(_1777_),
    .A(_1703_),
    .X(_1778_));
 sg13g2_nor3_1 _4114_ (.A(_1703_),
    .B(_1770_),
    .C(_1777_),
    .Y(_1779_));
 sg13g2_o21ai_1 _4115_ (.B1(_1754_),
    .Y(_1780_),
    .A1(_1768_),
    .A2(_1779_));
 sg13g2_or3_1 _4116_ (.A(_1754_),
    .B(_1768_),
    .C(_1779_),
    .X(_1781_));
 sg13g2_nand3_1 _4117_ (.B(_1780_),
    .C(_1781_),
    .A(_1236_),
    .Y(_1782_));
 sg13g2_nor2b_1 _4118_ (.A(_1778_),
    .B_N(_1782_),
    .Y(_1783_));
 sg13g2_nand4_1 _4119_ (.B(_1778_),
    .C(_1780_),
    .A(_1236_),
    .Y(_1784_),
    .D(_1781_));
 sg13g2_nand2_1 _4120_ (.Y(_1785_),
    .A(_1776_),
    .B(_1777_));
 sg13g2_o21ai_1 _4121_ (.B1(_1770_),
    .Y(_1786_),
    .A1(_1703_),
    .A2(_1777_));
 sg13g2_and2_1 _4122_ (.A(_1767_),
    .B(_1772_),
    .X(_1787_));
 sg13g2_nor3_1 _4123_ (.A(_1294_),
    .B(_1779_),
    .C(_1787_),
    .Y(_1788_));
 sg13g2_nand4_1 _4124_ (.B(_1785_),
    .C(_1786_),
    .A(_1784_),
    .Y(_1789_),
    .D(_1788_));
 sg13g2_o21ai_1 _4125_ (.B1(_1297_),
    .Y(_1790_),
    .A1(_1783_),
    .A2(_1789_));
 sg13g2_o21ai_1 _4126_ (.B1(_1592_),
    .Y(_1791_),
    .A1(_1398_),
    .A2(_1591_));
 sg13g2_a21o_1 _4127_ (.A2(_1591_),
    .A1(_1398_),
    .B1(_1791_),
    .X(_1792_));
 sg13g2_nand2_1 _4128_ (.Y(_0377_),
    .A(_1790_),
    .B(_1792_));
 sg13g2_nand2_1 _4129_ (.Y(_1793_),
    .A(_1495_),
    .B(_1694_));
 sg13g2_or2_1 _4130_ (.X(_1794_),
    .B(_1793_),
    .A(_1791_));
 sg13g2_nand3_1 _4131_ (.B(_1792_),
    .C(_1794_),
    .A(_1790_),
    .Y(_0376_));
 sg13g2_nand2_1 _4132_ (.Y(_1795_),
    .A(_1496_),
    .B(_1591_));
 sg13g2_or3_1 _4133_ (.A(_1398_),
    .B(_1591_),
    .C(_1700_),
    .X(_1796_));
 sg13g2_nand3_1 _4134_ (.B(_1795_),
    .C(_1796_),
    .A(_1592_),
    .Y(_1797_));
 sg13g2_nand2_2 _4135_ (.Y(_0378_),
    .A(_1790_),
    .B(_1797_));
 sg13g2_nand2b_1 _4136_ (.Y(_1798_),
    .B(_1697_),
    .A_N(_1594_));
 sg13g2_nand2b_1 _4137_ (.Y(_1799_),
    .B(_1694_),
    .A_N(_1798_));
 sg13g2_xor2_1 _4138_ (.B(_1012_),
    .A(_1011_),
    .X(_1800_));
 sg13g2_xor2_1 _4139_ (.B(_1757_),
    .A(_1011_),
    .X(_1801_));
 sg13g2_nand2_2 _4140_ (.Y(_1802_),
    .A(_1018_),
    .B(_1082_));
 sg13g2_nand3_1 _4141_ (.B(_1082_),
    .C(_1142_),
    .A(_1018_),
    .Y(_1803_));
 sg13g2_xnor2_1 _4142_ (.Y(_1804_),
    .A(_1718_),
    .B(_1802_));
 sg13g2_inv_1 _4143_ (.Y(_1805_),
    .A(_1804_));
 sg13g2_nand3_1 _4144_ (.B(_1082_),
    .C(_1121_),
    .A(_1018_),
    .Y(_1806_));
 sg13g2_xnor2_1 _4145_ (.Y(_1807_),
    .A(_1713_),
    .B(_1806_));
 sg13g2_inv_1 _4146_ (.Y(_1808_),
    .A(_1807_));
 sg13g2_nor2_2 _4147_ (.A(_1160_),
    .B(_1806_),
    .Y(_1809_));
 sg13g2_xor2_1 _4148_ (.B(_1809_),
    .A(_1723_),
    .X(_1810_));
 sg13g2_xnor2_1 _4149_ (.Y(_1811_),
    .A(_1723_),
    .B(_1809_));
 sg13g2_nor2_1 _4150_ (.A(_1807_),
    .B(_1811_),
    .Y(_1812_));
 sg13g2_xor2_1 _4151_ (.B(_1803_),
    .A(_1717_),
    .X(_1813_));
 sg13g2_nand3_1 _4152_ (.B(_1810_),
    .C(_1813_),
    .A(_1808_),
    .Y(_1814_));
 sg13g2_nor2b_1 _4153_ (.A(_1812_),
    .B_N(_1813_),
    .Y(_1815_));
 sg13g2_o21ai_1 _4154_ (.B1(_1813_),
    .Y(_1816_),
    .A1(_1807_),
    .A2(_1811_));
 sg13g2_nand4_1 _4155_ (.B(_1808_),
    .C(_1811_),
    .A(_1804_),
    .Y(_1817_),
    .D(_1813_));
 sg13g2_a221oi_1 _4156_ (.B2(_1811_),
    .C1(_1805_),
    .B1(_1817_),
    .A1(_1812_),
    .Y(_1818_),
    .A2(_1813_));
 sg13g2_a21oi_1 _4157_ (.A1(_1810_),
    .A2(_1814_),
    .Y(_1819_),
    .B1(_1804_));
 sg13g2_or2_1 _4158_ (.X(_1820_),
    .B(_1819_),
    .A(_1818_));
 sg13g2_xor2_1 _4159_ (.B(_1729_),
    .A(_1018_),
    .X(_1821_));
 sg13g2_nor4_1 _4160_ (.A(_1816_),
    .B(_1818_),
    .C(_1819_),
    .D(_1821_),
    .Y(_1822_));
 sg13g2_or3_1 _4161_ (.A(_1816_),
    .B(_1820_),
    .C(_1821_),
    .X(_1823_));
 sg13g2_a21oi_1 _4162_ (.A1(_1810_),
    .A2(_1813_),
    .Y(_1824_),
    .B1(_1807_));
 sg13g2_a21o_1 _4163_ (.A2(_1818_),
    .A1(_1815_),
    .B1(_1824_),
    .X(_1825_));
 sg13g2_a21oi_1 _4164_ (.A1(_1817_),
    .A2(_1825_),
    .Y(_1826_),
    .B1(_1822_));
 sg13g2_xnor2_1 _4165_ (.Y(_1827_),
    .A(_1821_),
    .B(_1826_));
 sg13g2_xnor2_1 _4166_ (.Y(_1828_),
    .A(_1009_),
    .B(_1017_));
 sg13g2_xnor2_1 _4167_ (.Y(_1829_),
    .A(_1073_),
    .B(_1706_));
 sg13g2_xor2_1 _4168_ (.B(_1829_),
    .A(_1828_),
    .X(_1830_));
 sg13g2_nor3_1 _4169_ (.A(_1820_),
    .B(_1821_),
    .C(_1826_),
    .Y(_1831_));
 sg13g2_xnor2_1 _4170_ (.Y(_1832_),
    .A(_1816_),
    .B(_1818_));
 sg13g2_o21ai_1 _4171_ (.B1(_1823_),
    .Y(_1833_),
    .A1(_1831_),
    .A2(_1832_));
 sg13g2_or2_1 _4172_ (.X(_1834_),
    .B(_1830_),
    .A(_1827_));
 sg13g2_or3_1 _4173_ (.A(_1820_),
    .B(_1827_),
    .C(_1830_),
    .X(_1835_));
 sg13g2_nand2_1 _4174_ (.Y(_1836_),
    .A(_1830_),
    .B(_1833_));
 sg13g2_a21o_1 _4175_ (.A2(_1835_),
    .A1(_1833_),
    .B1(_1830_),
    .X(_1837_));
 sg13g2_xor2_1 _4176_ (.B(_1016_),
    .A(_1013_),
    .X(_1838_));
 sg13g2_xnor2_1 _4177_ (.Y(_1839_),
    .A(_0995_),
    .B(_1192_));
 sg13g2_xnor2_1 _4178_ (.Y(_1840_),
    .A(_1838_),
    .B(_1839_));
 sg13g2_o21ai_1 _4179_ (.B1(_1820_),
    .Y(_1841_),
    .A1(_1821_),
    .A2(_1826_));
 sg13g2_nand2b_1 _4180_ (.Y(_1842_),
    .B(_1841_),
    .A_N(_1831_));
 sg13g2_inv_1 _4181_ (.Y(_1843_),
    .A(_1842_));
 sg13g2_a21oi_1 _4182_ (.A1(_1820_),
    .A2(_1833_),
    .Y(_1844_),
    .B1(_1834_));
 sg13g2_o21ai_1 _4183_ (.B1(_1835_),
    .Y(_1845_),
    .A1(_1843_),
    .A2(_1844_));
 sg13g2_and2_1 _4184_ (.A(_1836_),
    .B(_1837_),
    .X(_1846_));
 sg13g2_inv_1 _4185_ (.Y(_1847_),
    .A(_1846_));
 sg13g2_nand3b_1 _4186_ (.B(_1836_),
    .C(_1837_),
    .Y(_1848_),
    .A_N(_1827_));
 sg13g2_a21o_2 _4187_ (.A2(_1848_),
    .A1(_1845_),
    .B1(_1840_),
    .X(_1849_));
 sg13g2_o21ai_1 _4188_ (.B1(_1837_),
    .Y(_1850_),
    .A1(_1847_),
    .A2(_1849_));
 sg13g2_xnor2_1 _4189_ (.Y(_1851_),
    .A(_1827_),
    .B(_1850_));
 sg13g2_nand2_1 _4190_ (.Y(_1852_),
    .A(_1840_),
    .B(_1845_));
 sg13g2_nand2_2 _4191_ (.Y(_1853_),
    .A(_1849_),
    .B(_1852_));
 sg13g2_nor2_1 _4192_ (.A(_1847_),
    .B(_1853_),
    .Y(_1854_));
 sg13g2_o21ai_1 _4193_ (.B1(_1801_),
    .Y(_1855_),
    .A1(_1851_),
    .A2(_1854_));
 sg13g2_or2_1 _4194_ (.X(_1856_),
    .B(_1851_),
    .A(_1801_));
 sg13g2_and2_1 _4195_ (.A(_1855_),
    .B(_1856_),
    .X(_1857_));
 sg13g2_mux2_1 _4196_ (.A0(_1005_),
    .A1(_1060_),
    .S(_1010_),
    .X(_1858_));
 sg13g2_xnor2_1 _4197_ (.Y(_1859_),
    .A(_1702_),
    .B(_1858_));
 sg13g2_inv_1 _4198_ (.Y(_1860_),
    .A(_1859_));
 sg13g2_nand3_1 _4199_ (.B(_1856_),
    .C(_1859_),
    .A(_1855_),
    .Y(_1861_));
 sg13g2_or2_1 _4200_ (.X(_1862_),
    .B(_1861_),
    .A(_1853_));
 sg13g2_o21ai_1 _4201_ (.B1(_1849_),
    .Y(_1863_),
    .A1(_1853_),
    .A2(_1855_));
 sg13g2_xnor2_1 _4202_ (.Y(_1864_),
    .A(_1846_),
    .B(_1863_));
 sg13g2_a21o_1 _4203_ (.A2(_1864_),
    .A1(_1862_),
    .B1(_1860_),
    .X(_1865_));
 sg13g2_a21oi_1 _4204_ (.A1(_1853_),
    .A2(_1864_),
    .Y(_1866_),
    .B1(_1861_));
 sg13g2_xor2_1 _4205_ (.B(_1855_),
    .A(_1853_),
    .X(_1867_));
 sg13g2_o21ai_1 _4206_ (.B1(_1862_),
    .Y(_1868_),
    .A1(_1866_),
    .A2(_1867_));
 sg13g2_nor2b_2 _4207_ (.A(_0994_),
    .B_N(_1059_),
    .Y(_1869_));
 sg13g2_nand2_2 _4208_ (.Y(_1870_),
    .A(_1192_),
    .B(_1869_));
 sg13g2_xor2_1 _4209_ (.B(_1869_),
    .A(_1192_),
    .X(_1871_));
 sg13g2_xnor2_1 _4210_ (.Y(_1872_),
    .A(_1838_),
    .B(_1871_));
 sg13g2_inv_1 _4211_ (.Y(_1873_),
    .A(_1872_));
 sg13g2_nor2_1 _4212_ (.A(_1073_),
    .B(_1870_),
    .Y(_1874_));
 sg13g2_xnor2_1 _4213_ (.Y(_1875_),
    .A(_1018_),
    .B(_1874_));
 sg13g2_nor4_2 _4214_ (.A(_1073_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1876_),
    .D(_1870_));
 sg13g2_xnor2_1 _4215_ (.Y(_1877_),
    .A(_1089_),
    .B(_1875_));
 sg13g2_nand2_1 _4216_ (.Y(_1878_),
    .A(_1145_),
    .B(_1876_));
 sg13g2_nand4_1 _4217_ (.B(_1154_),
    .C(_1155_),
    .A(_1145_),
    .Y(_1879_),
    .D(_1876_));
 sg13g2_xnor2_1 _4218_ (.Y(_1880_),
    .A(_1806_),
    .B(_1879_));
 sg13g2_xnor2_1 _4219_ (.Y(_1881_),
    .A(_1166_),
    .B(_1880_));
 sg13g2_a21oi_1 _4220_ (.A1(_1161_),
    .A2(_1162_),
    .Y(_1882_),
    .B1(_1879_));
 sg13g2_xnor2_1 _4221_ (.Y(_1883_),
    .A(_1809_),
    .B(_1882_));
 sg13g2_xnor2_1 _4222_ (.Y(_1884_),
    .A(_1139_),
    .B(_1883_));
 sg13g2_xor2_1 _4223_ (.B(_1876_),
    .A(_1802_),
    .X(_1885_));
 sg13g2_xnor2_1 _4224_ (.Y(_1886_),
    .A(_1147_),
    .B(_1885_));
 sg13g2_xnor2_1 _4225_ (.Y(_1887_),
    .A(_1803_),
    .B(_1878_));
 sg13g2_xnor2_1 _4226_ (.Y(_1888_),
    .A(_1158_),
    .B(_1887_));
 sg13g2_nand3_1 _4227_ (.B(_1886_),
    .C(_1888_),
    .A(_1884_),
    .Y(_1889_));
 sg13g2_and2_1 _4228_ (.A(_1881_),
    .B(_1889_),
    .X(_1890_));
 sg13g2_nand3b_1 _4229_ (.B(_1886_),
    .C(_1888_),
    .Y(_1891_),
    .A_N(_1881_));
 sg13g2_nand3_1 _4230_ (.B(_1886_),
    .C(_1891_),
    .A(_1884_),
    .Y(_1892_));
 sg13g2_or2_1 _4231_ (.X(_1893_),
    .B(_1886_),
    .A(_1884_));
 sg13g2_nand2_1 _4232_ (.Y(_1894_),
    .A(_1892_),
    .B(_1893_));
 sg13g2_nor2b_1 _4233_ (.A(_1877_),
    .B_N(_1888_),
    .Y(_1895_));
 sg13g2_nand3_1 _4234_ (.B(_1893_),
    .C(_1895_),
    .A(_1892_),
    .Y(_1896_));
 sg13g2_nor2_1 _4235_ (.A(_1881_),
    .B(_1889_),
    .Y(_1897_));
 sg13g2_a21oi_2 _4236_ (.B1(_1897_),
    .Y(_1898_),
    .A2(_1896_),
    .A1(_1890_));
 sg13g2_xor2_1 _4237_ (.B(_1898_),
    .A(_1877_),
    .X(_1899_));
 sg13g2_xnor2_1 _4238_ (.Y(_1900_),
    .A(_1877_),
    .B(_1898_));
 sg13g2_xnor2_1 _4239_ (.Y(_1901_),
    .A(_1073_),
    .B(_1870_));
 sg13g2_xnor2_1 _4240_ (.Y(_1902_),
    .A(_1828_),
    .B(_1901_));
 sg13g2_nand2b_1 _4241_ (.Y(_1903_),
    .B(_1899_),
    .A_N(_1902_));
 sg13g2_or3_1 _4242_ (.A(_1894_),
    .B(_1900_),
    .C(_1902_),
    .X(_1904_));
 sg13g2_nor3_1 _4243_ (.A(_1877_),
    .B(_1894_),
    .C(_1898_),
    .Y(_1905_));
 sg13g2_xnor2_1 _4244_ (.Y(_1906_),
    .A(_1888_),
    .B(_1892_));
 sg13g2_xnor2_1 _4245_ (.Y(_1907_),
    .A(_1905_),
    .B(_1906_));
 sg13g2_a21oi_1 _4246_ (.A1(_1896_),
    .A2(_1897_),
    .Y(_1908_),
    .B1(_1890_));
 sg13g2_a21oi_1 _4247_ (.A1(_1890_),
    .A2(_1896_),
    .Y(_1909_),
    .B1(_1908_));
 sg13g2_a21oi_2 _4248_ (.B1(_1909_),
    .Y(_1910_),
    .A2(_1907_),
    .A1(_1904_));
 sg13g2_a21oi_1 _4249_ (.A1(_1904_),
    .A2(_1909_),
    .Y(_1911_),
    .B1(_1907_));
 sg13g2_a21oi_1 _4250_ (.A1(_1904_),
    .A2(_1907_),
    .Y(_1912_),
    .B1(_1911_));
 sg13g2_xor2_1 _4251_ (.B(_1910_),
    .A(_1902_),
    .X(_1913_));
 sg13g2_inv_1 _4252_ (.Y(_1914_),
    .A(_1913_));
 sg13g2_nor2_1 _4253_ (.A(_1872_),
    .B(_1900_),
    .Y(_1915_));
 sg13g2_nand2_1 _4254_ (.Y(_1916_),
    .A(_1913_),
    .B(_1915_));
 sg13g2_o21ai_1 _4255_ (.B1(_1894_),
    .Y(_1917_),
    .A1(_1877_),
    .A2(_1898_));
 sg13g2_nand2b_1 _4256_ (.Y(_1918_),
    .B(_1917_),
    .A_N(_1905_));
 sg13g2_o21ai_1 _4257_ (.B1(_1918_),
    .Y(_1919_),
    .A1(_1903_),
    .A2(_1910_));
 sg13g2_or3_1 _4258_ (.A(_1903_),
    .B(_1910_),
    .C(_1918_),
    .X(_1920_));
 sg13g2_nand2_1 _4259_ (.Y(_1921_),
    .A(_1919_),
    .B(_1920_));
 sg13g2_a22oi_1 _4260_ (.Y(_1922_),
    .B1(_1919_),
    .B2(_1920_),
    .A2(_1915_),
    .A1(_1913_));
 sg13g2_o21ai_1 _4261_ (.B1(_1873_),
    .Y(_1923_),
    .A1(_1912_),
    .A2(_1922_));
 sg13g2_or3_1 _4262_ (.A(_1873_),
    .B(_1912_),
    .C(_1921_),
    .X(_1924_));
 sg13g2_and2_1 _4263_ (.A(_1923_),
    .B(_1924_),
    .X(_1925_));
 sg13g2_inv_1 _4264_ (.Y(_1926_),
    .A(_1925_));
 sg13g2_xnor2_1 _4265_ (.Y(_1927_),
    .A(_0994_),
    .B(_1059_));
 sg13g2_or2_1 _4266_ (.X(_1928_),
    .B(_1927_),
    .A(_1800_));
 sg13g2_nand2_1 _4267_ (.Y(_1929_),
    .A(_1800_),
    .B(_1927_));
 sg13g2_nand2_1 _4268_ (.Y(_1930_),
    .A(_1928_),
    .B(_1929_));
 sg13g2_and4_1 _4269_ (.A(_1913_),
    .B(_1923_),
    .C(_1924_),
    .D(_1930_),
    .X(_1931_));
 sg13g2_o21ai_1 _4270_ (.B1(_1900_),
    .Y(_1932_),
    .A1(_1902_),
    .A2(_1910_));
 sg13g2_o21ai_1 _4271_ (.B1(_1932_),
    .Y(_1933_),
    .A1(_1903_),
    .A2(_1910_));
 sg13g2_nand4_1 _4272_ (.B(_1899_),
    .C(_1912_),
    .A(_1873_),
    .Y(_1934_),
    .D(_1913_));
 sg13g2_o21ai_1 _4273_ (.B1(_1933_),
    .Y(_1935_),
    .A1(_1914_),
    .A2(_1923_));
 sg13g2_nand2_1 _4274_ (.Y(_1936_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_a21oi_1 _4275_ (.A1(_1934_),
    .A2(_1935_),
    .Y(_1937_),
    .B1(_1931_));
 sg13g2_a21o_1 _4276_ (.A2(_1935_),
    .A1(_1934_),
    .B1(_1931_),
    .X(_1938_));
 sg13g2_a21oi_1 _4277_ (.A1(_1912_),
    .A2(_1916_),
    .Y(_1939_),
    .B1(_1921_));
 sg13g2_or2_1 _4278_ (.X(_1940_),
    .B(_1939_),
    .A(_1922_));
 sg13g2_inv_1 _4279_ (.Y(_1941_),
    .A(_1940_));
 sg13g2_nand4_1 _4280_ (.B(_1929_),
    .C(_1938_),
    .A(_1928_),
    .Y(_1942_),
    .D(_1940_));
 sg13g2_o21ai_1 _4281_ (.B1(_1930_),
    .Y(_1943_),
    .A1(_1937_),
    .A2(_1941_));
 sg13g2_xnor2_1 _4282_ (.Y(_1944_),
    .A(_1059_),
    .B(_1858_));
 sg13g2_inv_1 _4283_ (.Y(_1945_),
    .A(_1944_));
 sg13g2_nor2_1 _4284_ (.A(_1931_),
    .B(_1940_),
    .Y(_1946_));
 sg13g2_nor2_1 _4285_ (.A(_1936_),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_nor2_1 _4286_ (.A(_1937_),
    .B(_1947_),
    .Y(_1948_));
 sg13g2_nand2_1 _4287_ (.Y(_1949_),
    .A(_1942_),
    .B(_1943_));
 sg13g2_nand4_1 _4288_ (.B(_1942_),
    .C(_1943_),
    .A(_1925_),
    .Y(_1950_),
    .D(_1945_));
 sg13g2_xnor2_1 _4289_ (.Y(_1951_),
    .A(_1913_),
    .B(_1923_));
 sg13g2_a221oi_1 _4290_ (.B2(_1940_),
    .C1(_1926_),
    .B1(_1938_),
    .A1(_1928_),
    .Y(_1952_),
    .A2(_1929_));
 sg13g2_xnor2_1 _4291_ (.Y(_1953_),
    .A(_1951_),
    .B(_1952_));
 sg13g2_a21oi_1 _4292_ (.A1(_1950_),
    .A2(_1953_),
    .Y(_1954_),
    .B1(_1948_));
 sg13g2_or2_1 _4293_ (.X(_1955_),
    .B(_1954_),
    .A(_1944_));
 sg13g2_o21ai_1 _4294_ (.B1(_1943_),
    .Y(_1956_),
    .A1(_1944_),
    .A2(_1954_));
 sg13g2_and3_1 _4295_ (.X(_1957_),
    .A(_1925_),
    .B(_1942_),
    .C(_1956_));
 sg13g2_a21oi_1 _4296_ (.A1(_1942_),
    .A2(_1956_),
    .Y(_1958_),
    .B1(_1925_));
 sg13g2_nand2_1 _4297_ (.Y(_1959_),
    .A(_1944_),
    .B(_1954_));
 sg13g2_and4_1 _4298_ (.A(_1942_),
    .B(_1943_),
    .C(_1955_),
    .D(_1959_),
    .X(_1960_));
 sg13g2_inv_1 _4299_ (.Y(_1961_),
    .A(_1960_));
 sg13g2_o21ai_1 _4300_ (.B1(_1960_),
    .Y(_1962_),
    .A1(_1957_),
    .A2(_1958_));
 sg13g2_a21o_2 _4301_ (.A2(_1962_),
    .A1(_1868_),
    .B1(_1235_),
    .X(_1963_));
 sg13g2_and2_1 _4302_ (.A(_1860_),
    .B(_1864_),
    .X(_1964_));
 sg13g2_a21o_1 _4303_ (.A2(_1865_),
    .A1(_1235_),
    .B1(_1964_),
    .X(_1965_));
 sg13g2_o21ai_1 _4304_ (.B1(_1236_),
    .Y(_1966_),
    .A1(_1957_),
    .A2(_1958_));
 sg13g2_a21oi_1 _4305_ (.A1(_1860_),
    .A2(_1864_),
    .Y(_1967_),
    .B1(_1857_));
 sg13g2_xnor2_1 _4306_ (.Y(_1968_),
    .A(_1949_),
    .B(_1955_));
 sg13g2_mux2_1 _4307_ (.A0(_1953_),
    .A1(_1948_),
    .S(_1950_),
    .X(_1969_));
 sg13g2_or4_1 _4308_ (.A(_0662_),
    .B(_1967_),
    .C(_1968_),
    .D(_1969_),
    .X(_1970_));
 sg13g2_a221oi_1 _4309_ (.B2(_1961_),
    .C1(_1970_),
    .B1(_1966_),
    .A1(_1857_),
    .Y(_1971_),
    .A2(_1965_));
 sg13g2_nand2_1 _4310_ (.Y(_1972_),
    .A(_1963_),
    .B(_1971_));
 sg13g2_nand2_1 _4311_ (.Y(_1973_),
    .A(_0662_),
    .B(_1591_));
 sg13g2_a21oi_1 _4312_ (.A1(_1398_),
    .A2(_1700_),
    .Y(_1974_),
    .B1(_1973_));
 sg13g2_nor2b_1 _4313_ (.A(_1697_),
    .B_N(_1974_),
    .Y(_1975_));
 sg13g2_a21oi_2 _4314_ (.B1(_1975_),
    .Y(_1976_),
    .A2(_1971_),
    .A1(_1963_));
 sg13g2_nor2_1 _4315_ (.A(net747),
    .B(_1976_),
    .Y(_0381_));
 sg13g2_o21ai_1 _4316_ (.B1(_1799_),
    .Y(_0379_),
    .A1(net747),
    .A2(_1976_));
 sg13g2_o21ai_1 _4317_ (.B1(_1798_),
    .Y(_0380_),
    .A1(net747),
    .A2(_1976_));
 sg13g2_nand3_1 _4318_ (.B(_1699_),
    .C(_1793_),
    .A(_1399_),
    .Y(_1977_));
 sg13g2_a22oi_1 _4319_ (.Y(_1978_),
    .B1(_1974_),
    .B2(_1977_),
    .A2(_1698_),
    .A1(_1593_));
 sg13g2_a21oi_1 _4320_ (.A1(_1972_),
    .A2(_1978_),
    .Y(_0382_),
    .B1(net747));
 sg13g2_nand3_1 _4321_ (.B(_1693_),
    .C(_1974_),
    .A(net797),
    .Y(_1979_));
 sg13g2_and2_1 _4322_ (.A(_1799_),
    .B(_1979_),
    .X(_1980_));
 sg13g2_o21ai_1 _4323_ (.B1(_1980_),
    .Y(_0383_),
    .A1(net748),
    .A2(_1976_));
 sg13g2_xnor2_1 _4324_ (.Y(_1981_),
    .A(\tmds_red.n102 ),
    .B(_0914_));
 sg13g2_a21oi_1 _4325_ (.A1(net606),
    .A2(_1981_),
    .Y(_0384_),
    .B1(net747));
 sg13g2_xor2_1 _4326_ (.B(_0882_),
    .A(\tmds_red.n114 ),
    .X(_1982_));
 sg13g2_o21ai_1 _4327_ (.B1(net606),
    .Y(_1983_),
    .A1(_0914_),
    .A2(_1982_));
 sg13g2_a21oi_1 _4328_ (.A1(_0914_),
    .A2(_1982_),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_nor2_1 _4329_ (.A(net747),
    .B(_1984_),
    .Y(_0385_));
 sg13g2_xnor2_1 _4330_ (.Y(_1985_),
    .A(\tmds_red.n126 ),
    .B(_0882_));
 sg13g2_xnor2_1 _4331_ (.Y(_1986_),
    .A(_0910_),
    .B(_1985_));
 sg13g2_xor2_1 _4332_ (.B(_1985_),
    .A(net547),
    .X(_1987_));
 sg13g2_o21ai_1 _4333_ (.B1(net606),
    .Y(_1988_),
    .A1(_0906_),
    .A2(_1987_));
 sg13g2_a21oi_1 _4334_ (.A1(_0906_),
    .A2(_1986_),
    .Y(_1989_),
    .B1(_1988_));
 sg13g2_nor2_1 _4335_ (.A(net747),
    .B(_1989_),
    .Y(_0386_));
 sg13g2_nor2b_1 _4336_ (.A(net547),
    .B_N(net607),
    .Y(_1990_));
 sg13g2_nor2_1 _4337_ (.A(net749),
    .B(_1990_),
    .Y(_0387_));
 sg13g2_nor2b_1 _4338_ (.A(_0914_),
    .B_N(net606),
    .Y(_1991_));
 sg13g2_nor2_1 _4339_ (.A(net747),
    .B(_1991_),
    .Y(_0388_));
 sg13g2_a21oi_1 _4340_ (.A1(_0654_),
    .A2(net606),
    .Y(_0505_),
    .B1(net748));
 sg13g2_o21ai_1 _4341_ (.B1(net606),
    .Y(_1992_),
    .A1(\tmds_green.n126 ),
    .A2(_0860_));
 sg13g2_a21oi_1 _4342_ (.A1(_0860_),
    .A2(_0864_),
    .Y(_1993_),
    .B1(_1992_));
 sg13g2_nor2_1 _4343_ (.A(net748),
    .B(_1993_),
    .Y(_0506_));
 sg13g2_a21oi_1 _4344_ (.A1(\tmds_green.n100 ),
    .A2(net605),
    .Y(_0507_),
    .B1(net749));
 sg13g2_and2_1 _4345_ (.A(net606),
    .B(_0862_),
    .X(_1994_));
 sg13g2_a21oi_1 _4346_ (.A1(_0859_),
    .A2(_1994_),
    .Y(_0508_),
    .B1(net748));
 sg13g2_and2_1 _4347_ (.A(\tmds_red.dc_balancing_reg[0] ),
    .B(_0852_),
    .X(_0509_));
 sg13g2_xnor2_1 _4348_ (.Y(_1995_),
    .A(\tmds_red.n132 ),
    .B(\tmds_red.dc_balancing_reg[1] ));
 sg13g2_xnor2_1 _4349_ (.Y(_1996_),
    .A(\tmds_red.n114 ),
    .B(_1995_));
 sg13g2_xor2_1 _4350_ (.B(_1996_),
    .A(_0917_),
    .X(_1997_));
 sg13g2_nor2_1 _4351_ (.A(net571),
    .B(_1997_),
    .Y(_0510_));
 sg13g2_nand2_1 _4352_ (.Y(_1998_),
    .A(\tmds_red.dc_balancing_reg[2] ),
    .B(_0905_));
 sg13g2_xnor2_1 _4353_ (.Y(_1999_),
    .A(\tmds_red.dc_balancing_reg[2] ),
    .B(_0905_));
 sg13g2_inv_1 _4354_ (.Y(_2000_),
    .A(_1999_));
 sg13g2_nor2_1 _4355_ (.A(_0869_),
    .B(_0898_),
    .Y(_2001_));
 sg13g2_a21oi_1 _4356_ (.A1(_0665_),
    .A2(_0869_),
    .Y(_2002_),
    .B1(_2001_));
 sg13g2_inv_1 _4357_ (.Y(_2003_),
    .A(_2002_));
 sg13g2_xnor2_1 _4358_ (.Y(_2004_),
    .A(_1999_),
    .B(_2003_));
 sg13g2_or2_1 _4359_ (.X(_2005_),
    .B(_2004_),
    .A(_1996_));
 sg13g2_nor2_1 _4360_ (.A(net547),
    .B(_2005_),
    .Y(_2006_));
 sg13g2_inv_1 _4361_ (.Y(_2007_),
    .A(_2006_));
 sg13g2_xor2_1 _4362_ (.B(_2004_),
    .A(_1996_),
    .X(_2008_));
 sg13g2_o21ai_1 _4363_ (.B1(_2008_),
    .Y(_2009_),
    .A1(net548),
    .A2(_1996_));
 sg13g2_a21oi_1 _4364_ (.A1(_2007_),
    .A2(_2009_),
    .Y(_2010_),
    .B1(_0911_));
 sg13g2_a21o_1 _4365_ (.A2(_0869_),
    .A1(\tmds_red.dc_balancing_reg[1] ),
    .B1(_2001_),
    .X(_2011_));
 sg13g2_xor2_1 _4366_ (.B(_2011_),
    .A(_1999_),
    .X(_2012_));
 sg13g2_nor2_1 _4367_ (.A(_1996_),
    .B(_2012_),
    .Y(_2013_));
 sg13g2_xor2_1 _4368_ (.B(_2012_),
    .A(_1996_),
    .X(_2014_));
 sg13g2_nor2_1 _4369_ (.A(net548),
    .B(_0906_),
    .Y(_2015_));
 sg13g2_a22oi_1 _4370_ (.Y(_2016_),
    .B1(_2014_),
    .B2(_2015_),
    .A2(_2008_),
    .A1(_0913_));
 sg13g2_nand2_1 _4371_ (.Y(_2017_),
    .A(net548),
    .B(_1996_));
 sg13g2_nor2b_1 _4372_ (.A(_2014_),
    .B_N(_2017_),
    .Y(_2018_));
 sg13g2_nor2_1 _4373_ (.A(_2012_),
    .B(_2017_),
    .Y(_2019_));
 sg13g2_nor3_1 _4374_ (.A(_0910_),
    .B(_2018_),
    .C(_2019_),
    .Y(_2020_));
 sg13g2_nor2_1 _4375_ (.A(_2010_),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_a21oi_1 _4376_ (.A1(_2016_),
    .A2(_2021_),
    .Y(_0511_),
    .B1(net571));
 sg13g2_o21ai_1 _4377_ (.B1(_2005_),
    .Y(_2022_),
    .A1(_1999_),
    .A2(_2003_));
 sg13g2_o21ai_1 _4378_ (.B1(_0905_),
    .Y(_2023_),
    .A1(_0901_),
    .A2(_0902_));
 sg13g2_xnor2_1 _4379_ (.Y(_2024_),
    .A(_0666_),
    .B(_2023_));
 sg13g2_nand2_1 _4380_ (.Y(_2025_),
    .A(_0907_),
    .B(_1998_));
 sg13g2_and2_1 _4381_ (.A(_2024_),
    .B(_2025_),
    .X(_2026_));
 sg13g2_xor2_1 _4382_ (.B(_2025_),
    .A(_2024_),
    .X(_2027_));
 sg13g2_xor2_1 _4383_ (.B(_2027_),
    .A(_2022_),
    .X(_2028_));
 sg13g2_nand2_1 _4384_ (.Y(_2029_),
    .A(_2007_),
    .B(_2028_));
 sg13g2_and2_1 _4385_ (.A(_2006_),
    .B(_2027_),
    .X(_2030_));
 sg13g2_a21oi_1 _4386_ (.A1(_2000_),
    .A2(_2011_),
    .Y(_2031_),
    .B1(_2013_));
 sg13g2_o21ai_1 _4387_ (.B1(_1998_),
    .Y(_2032_),
    .A1(_0903_),
    .A2(_0905_));
 sg13g2_xor2_1 _4388_ (.B(_2032_),
    .A(_2024_),
    .X(_2033_));
 sg13g2_nor2b_1 _4389_ (.A(_2031_),
    .B_N(_2033_),
    .Y(_2034_));
 sg13g2_xnor2_1 _4390_ (.Y(_2035_),
    .A(_2031_),
    .B(_2033_));
 sg13g2_and2_1 _4391_ (.A(_2019_),
    .B(_2035_),
    .X(_2036_));
 sg13g2_a21oi_1 _4392_ (.A1(_2024_),
    .A2(_2032_),
    .Y(_2037_),
    .B1(_2034_));
 sg13g2_a21oi_1 _4393_ (.A1(_0666_),
    .A2(_2023_),
    .Y(_2038_),
    .B1(_0902_));
 sg13g2_xnor2_1 _4394_ (.Y(_2039_),
    .A(\tmds_red.dc_balancing_reg[4] ),
    .B(_2038_));
 sg13g2_xnor2_1 _4395_ (.Y(_2040_),
    .A(_2037_),
    .B(_2039_));
 sg13g2_inv_1 _4396_ (.Y(_2041_),
    .A(_2040_));
 sg13g2_xnor2_1 _4397_ (.Y(_2042_),
    .A(_2019_),
    .B(_2035_));
 sg13g2_nand2b_1 _4398_ (.Y(_2043_),
    .B(_2042_),
    .A_N(_0910_));
 sg13g2_nand3b_1 _4399_ (.B(_0910_),
    .C(_2029_),
    .Y(_2044_),
    .A_N(_2030_));
 sg13g2_nand3_1 _4400_ (.B(_2043_),
    .C(_2044_),
    .A(_0906_),
    .Y(_2045_));
 sg13g2_a22oi_1 _4401_ (.Y(_2046_),
    .B1(_2035_),
    .B2(_2015_),
    .A2(_2028_),
    .A1(_0913_));
 sg13g2_a21oi_1 _4402_ (.A1(_2045_),
    .A2(_2046_),
    .Y(_0512_),
    .B1(net571));
 sg13g2_nor3_1 _4403_ (.A(_0910_),
    .B(_2036_),
    .C(_2041_),
    .Y(_2047_));
 sg13g2_a21oi_1 _4404_ (.A1(_2022_),
    .A2(_2027_),
    .Y(_2048_),
    .B1(_2026_));
 sg13g2_a21oi_1 _4405_ (.A1(\tmds_red.dc_balancing_reg[3] ),
    .A2(_2023_),
    .Y(_2049_),
    .B1(_0902_));
 sg13g2_xnor2_1 _4406_ (.Y(_2050_),
    .A(_0664_),
    .B(_2049_));
 sg13g2_xnor2_1 _4407_ (.Y(_2051_),
    .A(_2048_),
    .B(_2050_));
 sg13g2_o21ai_1 _4408_ (.B1(_0910_),
    .Y(_2052_),
    .A1(_2030_),
    .A2(_2051_));
 sg13g2_a21oi_1 _4409_ (.A1(_2030_),
    .A2(_2051_),
    .Y(_2053_),
    .B1(_2052_));
 sg13g2_o21ai_1 _4410_ (.B1(_0906_),
    .Y(_2054_),
    .A1(_2047_),
    .A2(_2053_));
 sg13g2_a22oi_1 _4411_ (.Y(_2055_),
    .B1(_2051_),
    .B2(_0913_),
    .A2(_2040_),
    .A1(_2015_));
 sg13g2_a21oi_1 _4412_ (.A1(_2054_),
    .A2(_2055_),
    .Y(_0513_),
    .B1(net572));
 sg13g2_or4_1 _4413_ (.A(\tmds_blue.dc_balancing_reg[0] ),
    .B(\tmds_blue.dc_balancing_reg[1] ),
    .C(\tmds_blue.dc_balancing_reg[3] ),
    .D(\tmds_blue.dc_balancing_reg[2] ),
    .X(_2056_));
 sg13g2_nor2_2 _4414_ (.A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_2056_),
    .Y(_2057_));
 sg13g2_nand2b_1 _4415_ (.Y(_2058_),
    .B(\tmds_blue.dc_balancing_reg[4] ),
    .A_N(\tmds_blue.n193 ));
 sg13g2_nand3_1 _4416_ (.B(_0655_),
    .C(_2056_),
    .A(\tmds_blue.n193 ),
    .Y(_2059_));
 sg13g2_and2_1 _4417_ (.A(_2058_),
    .B(_2059_),
    .X(_2060_));
 sg13g2_nand2_2 _4418_ (.Y(_2061_),
    .A(_2058_),
    .B(_2059_));
 sg13g2_xnor2_1 _4419_ (.Y(_2062_),
    .A(net602),
    .B(_2060_));
 sg13g2_nand2b_2 _4420_ (.Y(_2063_),
    .B(_2062_),
    .A_N(_2057_));
 sg13g2_o21ai_1 _4421_ (.B1(net799),
    .Y(_2064_),
    .A1(net605),
    .A2(hsync));
 sg13g2_a21oi_1 _4422_ (.A1(net605),
    .A2(_2063_),
    .Y(_0610_),
    .B1(_2064_));
 sg13g2_nand2b_1 _4423_ (.Y(_2065_),
    .B(\tmds_blue.n193 ),
    .A_N(net603));
 sg13g2_xnor2_1 _4424_ (.Y(_2066_),
    .A(net604),
    .B(\tmds_blue.n193 ));
 sg13g2_o21ai_1 _4425_ (.B1(net605),
    .Y(_2067_),
    .A1(_2056_),
    .A2(_2066_));
 sg13g2_nor2_2 _4426_ (.A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_nor2_1 _4427_ (.A(_2064_),
    .B(_2068_),
    .Y(_0611_));
 sg13g2_o21ai_1 _4428_ (.B1(net799),
    .Y(_2069_),
    .A1(net605),
    .A2(_0667_));
 sg13g2_nor2_1 _4429_ (.A(_2068_),
    .B(_2069_),
    .Y(_0612_));
 sg13g2_a21oi_1 _4430_ (.A1(net603),
    .A2(_2057_),
    .Y(_2070_),
    .B1(_2061_));
 sg13g2_xnor2_1 _4431_ (.Y(_2071_),
    .A(\tmds_blue.n126 ),
    .B(_2066_));
 sg13g2_xor2_1 _4432_ (.B(_2071_),
    .A(_2070_),
    .X(_2072_));
 sg13g2_a21oi_1 _4433_ (.A1(net605),
    .A2(_2072_),
    .Y(_0615_),
    .B1(_2069_));
 sg13g2_xnor2_1 _4434_ (.Y(_2073_),
    .A(net604),
    .B(\tmds_blue.n132 ));
 sg13g2_xnor2_1 _4435_ (.Y(_2074_),
    .A(_2072_),
    .B(_2073_));
 sg13g2_a21oi_1 _4436_ (.A1(net605),
    .A2(_2074_),
    .Y(_0616_),
    .B1(_2064_));
 sg13g2_a21oi_1 _4437_ (.A1(net604),
    .A2(net605),
    .Y(_0617_),
    .B1(_2069_));
 sg13g2_xnor2_1 _4438_ (.Y(_2075_),
    .A(hsync),
    .B(\tmds_blue.vsync ));
 sg13g2_nand2_1 _4439_ (.Y(_2076_),
    .A(net801),
    .B(_2075_));
 sg13g2_a22oi_1 _4440_ (.Y(_0618_),
    .B1(_2076_),
    .B2(net572),
    .A2(_2070_),
    .A1(net607));
 sg13g2_nand2b_1 _4441_ (.Y(_2077_),
    .B(\tmds_green.dc_balancing_reg[1] ),
    .A_N(net599));
 sg13g2_nand2_1 _4442_ (.Y(_2078_),
    .A(net599),
    .B(_0652_));
 sg13g2_and3_2 _4443_ (.X(_2079_),
    .A(net600),
    .B(_2077_),
    .C(_2078_));
 sg13g2_a21oi_1 _4444_ (.A1(_2077_),
    .A2(_2078_),
    .Y(_2080_),
    .B1(net600));
 sg13g2_nor2_2 _4445_ (.A(_2079_),
    .B(_2080_),
    .Y(_2081_));
 sg13g2_o21ai_1 _4446_ (.B1(_0852_),
    .Y(_2082_),
    .A1(_0654_),
    .A2(_2081_));
 sg13g2_a21oi_1 _4447_ (.A1(_0654_),
    .A2(_2081_),
    .Y(_0619_),
    .B1(_2082_));
 sg13g2_nor2_1 _4448_ (.A(net599),
    .B(\tmds_green.n126 ),
    .Y(_2083_));
 sg13g2_nor3_1 _4449_ (.A(net600),
    .B(net599),
    .C(\tmds_green.n126 ),
    .Y(_2084_));
 sg13g2_nand2_1 _4450_ (.Y(_2085_),
    .A(net599),
    .B(\tmds_green.n126 ));
 sg13g2_nand3_1 _4451_ (.B(\tmds_green.n132 ),
    .C(\tmds_green.n126 ),
    .A(net600),
    .Y(_2086_));
 sg13g2_nor2_1 _4452_ (.A(net601),
    .B(_2083_),
    .Y(_2087_));
 sg13g2_nand2b_2 _4453_ (.Y(_2088_),
    .B(_2086_),
    .A_N(_2084_));
 sg13g2_nor2b_1 _4454_ (.A(\tmds_green.dc_balancing_reg[2] ),
    .B_N(_2088_),
    .Y(_2089_));
 sg13g2_xnor2_1 _4455_ (.Y(_2090_),
    .A(\tmds_green.dc_balancing_reg[2] ),
    .B(_2088_));
 sg13g2_o21ai_1 _4456_ (.B1(_0857_),
    .Y(_2091_),
    .A1(\tmds_green.dc_balancing_reg[1] ),
    .A2(_0858_));
 sg13g2_nor2_1 _4457_ (.A(_2090_),
    .B(_2091_),
    .Y(_2092_));
 sg13g2_nand2_1 _4458_ (.Y(_2093_),
    .A(_2090_),
    .B(_2091_));
 sg13g2_nand2b_1 _4459_ (.Y(_2094_),
    .B(_2093_),
    .A_N(_2092_));
 sg13g2_xor2_1 _4460_ (.B(_2094_),
    .A(_2079_),
    .X(_2095_));
 sg13g2_nand2b_1 _4461_ (.Y(_2096_),
    .B(_2090_),
    .A_N(_2078_));
 sg13g2_a21oi_2 _4462_ (.B1(_2090_),
    .Y(_2097_),
    .A2(_0652_),
    .A1(net599));
 sg13g2_nor2_1 _4463_ (.A(_0863_),
    .B(_2097_),
    .Y(_2098_));
 sg13g2_a22oi_1 _4464_ (.Y(_2099_),
    .B1(_2096_),
    .B2(_2098_),
    .A2(_2095_),
    .A1(_0863_));
 sg13g2_xnor2_1 _4465_ (.Y(_2100_),
    .A(_0860_),
    .B(_2099_));
 sg13g2_nor2_1 _4466_ (.A(net571),
    .B(_2100_),
    .Y(_0620_));
 sg13g2_xnor2_1 _4467_ (.Y(_2101_),
    .A(_0653_),
    .B(_2088_));
 sg13g2_inv_1 _4468_ (.Y(_2102_),
    .A(_2101_));
 sg13g2_a21o_1 _4469_ (.A2(_2085_),
    .A1(net600),
    .B1(_2089_),
    .X(_2103_));
 sg13g2_xnor2_1 _4470_ (.Y(_2104_),
    .A(_2102_),
    .B(_2103_));
 sg13g2_o21ai_1 _4471_ (.B1(_2093_),
    .Y(_2105_),
    .A1(_2081_),
    .A2(_2092_));
 sg13g2_nand2b_1 _4472_ (.Y(_2106_),
    .B(_2104_),
    .A_N(_2105_));
 sg13g2_xnor2_1 _4473_ (.Y(_2107_),
    .A(_2104_),
    .B(_2105_));
 sg13g2_nand3_1 _4474_ (.B(_2090_),
    .C(_2107_),
    .A(_2080_),
    .Y(_2108_));
 sg13g2_nand2_1 _4475_ (.Y(_2109_),
    .A(_0863_),
    .B(_2108_));
 sg13g2_a21oi_1 _4476_ (.A1(_2080_),
    .A2(_2090_),
    .Y(_2110_),
    .B1(_2107_));
 sg13g2_nor2_1 _4477_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_nor2_1 _4478_ (.A(_2087_),
    .B(_2089_),
    .Y(_2112_));
 sg13g2_inv_1 _4479_ (.Y(_2113_),
    .A(_2112_));
 sg13g2_xnor2_1 _4480_ (.Y(_2114_),
    .A(_2101_),
    .B(_2112_));
 sg13g2_xnor2_1 _4481_ (.Y(_2115_),
    .A(_2097_),
    .B(_2114_));
 sg13g2_nor2_1 _4482_ (.A(_0863_),
    .B(_2115_),
    .Y(_2116_));
 sg13g2_nor3_1 _4483_ (.A(_0856_),
    .B(_2111_),
    .C(_2116_),
    .Y(_2117_));
 sg13g2_nor2_1 _4484_ (.A(net571),
    .B(_2117_),
    .Y(_0621_));
 sg13g2_o21ai_1 _4485_ (.B1(_2106_),
    .Y(_2118_),
    .A1(_2101_),
    .A2(_2103_));
 sg13g2_a21oi_1 _4486_ (.A1(\tmds_green.dc_balancing_reg[3] ),
    .A2(_2086_),
    .Y(_2119_),
    .B1(_2084_));
 sg13g2_xnor2_1 _4487_ (.Y(_2120_),
    .A(_0654_),
    .B(_2119_));
 sg13g2_xnor2_1 _4488_ (.Y(_2121_),
    .A(_2118_),
    .B(_2120_));
 sg13g2_nor2_1 _4489_ (.A(_2109_),
    .B(_2121_),
    .Y(_2122_));
 sg13g2_nand2_1 _4490_ (.Y(_2123_),
    .A(_2077_),
    .B(_2090_));
 sg13g2_nand3_1 _4491_ (.B(_2114_),
    .C(_2123_),
    .A(net600),
    .Y(_2124_));
 sg13g2_or2_1 _4492_ (.X(_2125_),
    .B(_2124_),
    .A(_2097_));
 sg13g2_a221oi_1 _4493_ (.B2(net600),
    .C1(_2097_),
    .B1(_2123_),
    .A1(_2102_),
    .Y(_2126_),
    .A2(_2112_));
 sg13g2_a21oi_1 _4494_ (.A1(_2101_),
    .A2(_2113_),
    .Y(_2127_),
    .B1(_2126_));
 sg13g2_o21ai_1 _4495_ (.B1(_2086_),
    .Y(_2128_),
    .A1(_0653_),
    .A2(_2084_));
 sg13g2_xnor2_1 _4496_ (.Y(_2129_),
    .A(\tmds_green.dc_balancing_reg[4] ),
    .B(_2128_));
 sg13g2_xnor2_1 _4497_ (.Y(_2130_),
    .A(_2127_),
    .B(_2129_));
 sg13g2_a21oi_1 _4498_ (.A1(_2125_),
    .A2(_2130_),
    .Y(_2131_),
    .B1(_0863_));
 sg13g2_nor3_1 _4499_ (.A(_0856_),
    .B(_2122_),
    .C(_2131_),
    .Y(_2132_));
 sg13g2_nor2_1 _4500_ (.A(net572),
    .B(_2132_),
    .Y(_0622_));
 sg13g2_nor3_1 _4501_ (.A(net751),
    .B(\clockdiv.q0 ),
    .C(net406),
    .Y(_0623_));
 sg13g2_xnor2_1 _4502_ (.Y(_2133_),
    .A(\tmds_blue.n193 ),
    .B(\tmds_blue.dc_balancing_reg[1] ));
 sg13g2_xnor2_1 _4503_ (.Y(_2134_),
    .A(\tmds_blue.n132 ),
    .B(_2133_));
 sg13g2_xor2_1 _4504_ (.B(_2134_),
    .A(_2063_),
    .X(_2135_));
 sg13g2_nor2_1 _4505_ (.A(net572),
    .B(_2135_),
    .Y(_0624_));
 sg13g2_and2_1 _4506_ (.A(\tmds_blue.n126 ),
    .B(\tmds_blue.n132 ),
    .X(_2136_));
 sg13g2_nor3_1 _4507_ (.A(net603),
    .B(_2071_),
    .C(_2136_),
    .Y(_2137_));
 sg13g2_a21oi_1 _4508_ (.A1(_2065_),
    .A2(_2136_),
    .Y(_2138_),
    .B1(_2137_));
 sg13g2_xor2_1 _4509_ (.B(\tmds_blue.n193 ),
    .A(\tmds_blue.n132 ),
    .X(_2139_));
 sg13g2_nor2_2 _4510_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sg13g2_nand2b_1 _4511_ (.Y(_2141_),
    .B(_2140_),
    .A_N(\tmds_blue.dc_balancing_reg[2] ));
 sg13g2_xnor2_1 _4512_ (.Y(_2142_),
    .A(\tmds_blue.dc_balancing_reg[2] ),
    .B(_2140_));
 sg13g2_nand2b_1 _4513_ (.Y(_2143_),
    .B(_2139_),
    .A_N(_2138_));
 sg13g2_o21ai_1 _4514_ (.B1(_2143_),
    .Y(_2144_),
    .A1(\tmds_blue.dc_balancing_reg[1] ),
    .A2(_2139_));
 sg13g2_nor2_1 _4515_ (.A(_2142_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_xnor2_1 _4516_ (.Y(_2146_),
    .A(_2142_),
    .B(_2144_));
 sg13g2_nor2_1 _4517_ (.A(_2134_),
    .B(_2146_),
    .Y(_2147_));
 sg13g2_nand2_1 _4518_ (.Y(_2148_),
    .A(net602),
    .B(_2147_));
 sg13g2_xnor2_1 _4519_ (.Y(_2149_),
    .A(_2134_),
    .B(_2146_));
 sg13g2_o21ai_1 _4520_ (.B1(_2143_),
    .Y(_2150_),
    .A1(_0656_),
    .A2(_2139_));
 sg13g2_nand2b_1 _4521_ (.Y(_2151_),
    .B(_2150_),
    .A_N(_2142_));
 sg13g2_xnor2_1 _4522_ (.Y(_2152_),
    .A(_2142_),
    .B(_2150_));
 sg13g2_nand2b_1 _4523_ (.Y(_2153_),
    .B(_2152_),
    .A_N(_2134_));
 sg13g2_xor2_1 _4524_ (.B(_2152_),
    .A(_2134_),
    .X(_2154_));
 sg13g2_nand2_1 _4525_ (.Y(_2155_),
    .A(net602),
    .B(_2154_));
 sg13g2_nor2b_1 _4526_ (.A(net602),
    .B_N(_2152_),
    .Y(_2156_));
 sg13g2_nor2b_1 _4527_ (.A(_2134_),
    .B_N(net602),
    .Y(_2157_));
 sg13g2_o21ai_1 _4528_ (.B1(_2148_),
    .Y(_2158_),
    .A1(_2149_),
    .A2(_2157_));
 sg13g2_nor2_1 _4529_ (.A(_2060_),
    .B(_2156_),
    .Y(_2159_));
 sg13g2_a221oi_1 _4530_ (.B2(_2155_),
    .C1(_2057_),
    .B1(_2159_),
    .A1(_2060_),
    .Y(_2160_),
    .A2(_2158_));
 sg13g2_nand2b_1 _4531_ (.Y(_2161_),
    .B(_2149_),
    .A_N(net602));
 sg13g2_nand2_1 _4532_ (.Y(_2162_),
    .A(_2155_),
    .B(_2161_));
 sg13g2_a21oi_1 _4533_ (.A1(_2057_),
    .A2(_2162_),
    .Y(_2163_),
    .B1(net572));
 sg13g2_nor2b_1 _4534_ (.A(_2160_),
    .B_N(_2163_),
    .Y(_0625_));
 sg13g2_xnor2_1 _4535_ (.Y(_2164_),
    .A(\tmds_blue.dc_balancing_reg[3] ),
    .B(_2140_));
 sg13g2_nand2_1 _4536_ (.Y(_2165_),
    .A(net603),
    .B(_2136_));
 sg13g2_nand2_1 _4537_ (.Y(_2166_),
    .A(\tmds_blue.n193 ),
    .B(_2165_));
 sg13g2_nand2_1 _4538_ (.Y(_2167_),
    .A(_2141_),
    .B(_2166_));
 sg13g2_inv_1 _4539_ (.Y(_2168_),
    .A(_2167_));
 sg13g2_xor2_1 _4540_ (.B(_2167_),
    .A(_2164_),
    .X(_2169_));
 sg13g2_a21oi_1 _4541_ (.A1(_2151_),
    .A2(_2153_),
    .Y(_2170_),
    .B1(_2169_));
 sg13g2_a21oi_1 _4542_ (.A1(_2164_),
    .A2(_2168_),
    .Y(_2171_),
    .B1(_2170_));
 sg13g2_nand3_1 _4543_ (.B(\tmds_blue.n193 ),
    .C(_2136_),
    .A(net603),
    .Y(_2172_));
 sg13g2_o21ai_1 _4544_ (.B1(_2172_),
    .Y(_2173_),
    .A1(\tmds_blue.dc_balancing_reg[3] ),
    .A2(_2140_));
 sg13g2_xnor2_1 _4545_ (.Y(_2174_),
    .A(\tmds_blue.dc_balancing_reg[4] ),
    .B(_2173_));
 sg13g2_xnor2_1 _4546_ (.Y(_2175_),
    .A(_2171_),
    .B(_2174_));
 sg13g2_nor2_1 _4547_ (.A(_2145_),
    .B(_2147_),
    .Y(_2176_));
 sg13g2_o21ai_1 _4548_ (.B1(_2166_),
    .Y(_2177_),
    .A1(_2138_),
    .A2(_2139_));
 sg13g2_nand2_1 _4549_ (.Y(_2178_),
    .A(_2141_),
    .B(_2177_));
 sg13g2_nand3_1 _4550_ (.B(_2164_),
    .C(_2177_),
    .A(_2141_),
    .Y(_2179_));
 sg13g2_xor2_1 _4551_ (.B(_2178_),
    .A(_2164_),
    .X(_2180_));
 sg13g2_xor2_1 _4552_ (.B(_2180_),
    .A(_2176_),
    .X(_2181_));
 sg13g2_o21ai_1 _4553_ (.B1(_2057_),
    .Y(_2182_),
    .A1(net602),
    .A2(_2181_));
 sg13g2_a21oi_1 _4554_ (.A1(net602),
    .A2(_2175_),
    .Y(_2183_),
    .B1(_2182_));
 sg13g2_nor2_1 _4555_ (.A(_2148_),
    .B(_2181_),
    .Y(_2184_));
 sg13g2_inv_1 _4556_ (.Y(_2185_),
    .A(_2184_));
 sg13g2_nand3_1 _4557_ (.B(_2153_),
    .C(_2169_),
    .A(_2151_),
    .Y(_2186_));
 sg13g2_nor2b_1 _4558_ (.A(_2170_),
    .B_N(_2186_),
    .Y(_2187_));
 sg13g2_a21oi_1 _4559_ (.A1(_2134_),
    .A2(_2156_),
    .Y(_2188_),
    .B1(_2187_));
 sg13g2_nand3_1 _4560_ (.B(_2156_),
    .C(_2187_),
    .A(_2134_),
    .Y(_2189_));
 sg13g2_nand2b_1 _4561_ (.Y(_2190_),
    .B(_2189_),
    .A_N(_2188_));
 sg13g2_a21oi_1 _4562_ (.A1(_2148_),
    .A2(_2181_),
    .Y(_2191_),
    .B1(_2061_));
 sg13g2_a221oi_1 _4563_ (.B2(_2185_),
    .C1(_2057_),
    .B1(_2191_),
    .A1(_2061_),
    .Y(_2192_),
    .A2(_2190_));
 sg13g2_nor2_1 _4564_ (.A(_2183_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_nor2_1 _4565_ (.A(net572),
    .B(_2193_),
    .Y(_0626_));
 sg13g2_o21ai_1 _4566_ (.B1(_2179_),
    .Y(_2194_),
    .A1(_2176_),
    .A2(_2180_));
 sg13g2_o21ai_1 _4567_ (.B1(_2172_),
    .Y(_2195_),
    .A1(_0657_),
    .A2(_2140_));
 sg13g2_xnor2_1 _4568_ (.Y(_2196_),
    .A(_0655_),
    .B(_2195_));
 sg13g2_xnor2_1 _4569_ (.Y(_2197_),
    .A(_2194_),
    .B(_2196_));
 sg13g2_o21ai_1 _4570_ (.B1(_2060_),
    .Y(_2198_),
    .A1(_2184_),
    .A2(_2197_));
 sg13g2_nand3b_1 _4571_ (.B(_2189_),
    .C(_2061_),
    .Y(_2199_),
    .A_N(_2175_));
 sg13g2_a21oi_1 _4572_ (.A1(_2198_),
    .A2(_2199_),
    .Y(_2200_),
    .B1(_2057_));
 sg13g2_nor2_1 _4573_ (.A(_2183_),
    .B(_2200_),
    .Y(_2201_));
 sg13g2_nor2_1 _4574_ (.A(net572),
    .B(_2201_),
    .Y(_0627_));
 sg13g2_nor2_1 _4575_ (.A(net674),
    .B(net726),
    .Y(_0007_));
 sg13g2_nor2_1 _4576_ (.A(net674),
    .B(net726),
    .Y(_0008_));
 sg13g2_nor2_1 _4577_ (.A(net677),
    .B(net729),
    .Y(_0009_));
 sg13g2_nor2_1 _4578_ (.A(_0654_),
    .B(net571),
    .Y(_0272_));
 sg13g2_a21oi_1 _4579_ (.A1(_0882_),
    .A2(_0917_),
    .Y(_0277_),
    .B1(_0918_));
 sg13g2_nor2_1 _4580_ (.A(net665),
    .B(net717),
    .Y(_0010_));
 sg13g2_nor2_1 _4581_ (.A(net666),
    .B(net718),
    .Y(_0011_));
 sg13g2_nor2_1 _4582_ (.A(net665),
    .B(net717),
    .Y(_0012_));
 sg13g2_nor2_1 _4583_ (.A(net665),
    .B(net717),
    .Y(_0013_));
 sg13g2_nor2_1 _4584_ (.A(net652),
    .B(net704),
    .Y(_0014_));
 sg13g2_nor2_1 _4585_ (.A(net652),
    .B(net704),
    .Y(_0015_));
 sg13g2_nor2_1 _4586_ (.A(net657),
    .B(net709),
    .Y(_0016_));
 sg13g2_nor2_1 _4587_ (.A(net657),
    .B(net709),
    .Y(_0017_));
 sg13g2_nor2_1 _4588_ (.A(net685),
    .B(net737),
    .Y(_0018_));
 sg13g2_nor2_1 _4589_ (.A(net685),
    .B(net737),
    .Y(_0019_));
 sg13g2_nor2_1 _4590_ (.A(net686),
    .B(net738),
    .Y(_0020_));
 sg13g2_nor2_1 _4591_ (.A(net684),
    .B(net736),
    .Y(_0021_));
 sg13g2_nor2_1 _4592_ (.A(net649),
    .B(net701),
    .Y(_0022_));
 sg13g2_nor2_1 _4593_ (.A(net649),
    .B(net701),
    .Y(_0023_));
 sg13g2_nor2_1 _4594_ (.A(net649),
    .B(net701),
    .Y(_0024_));
 sg13g2_nor2_1 _4595_ (.A(net649),
    .B(net703),
    .Y(_0025_));
 sg13g2_nor2_1 _4596_ (.A(net665),
    .B(net717),
    .Y(_0026_));
 sg13g2_nor2_1 _4597_ (.A(net661),
    .B(net713),
    .Y(_0027_));
 sg13g2_nor2_1 _4598_ (.A(net662),
    .B(net714),
    .Y(_0028_));
 sg13g2_nor2_1 _4599_ (.A(net661),
    .B(net713),
    .Y(_0029_));
 sg13g2_nor2_1 _4600_ (.A(net660),
    .B(net712),
    .Y(_0030_));
 sg13g2_nor2_1 _4601_ (.A(net660),
    .B(net712),
    .Y(_0031_));
 sg13g2_nor2_1 _4602_ (.A(net662),
    .B(net714),
    .Y(_0032_));
 sg13g2_nor2_1 _4603_ (.A(net660),
    .B(net712),
    .Y(_0033_));
 sg13g2_nor2_1 _4604_ (.A(net683),
    .B(net734),
    .Y(_0034_));
 sg13g2_nor2_1 _4605_ (.A(net668),
    .B(net719),
    .Y(_0035_));
 sg13g2_nor2_1 _4606_ (.A(net684),
    .B(net736),
    .Y(_0036_));
 sg13g2_nor2_1 _4607_ (.A(net683),
    .B(net719),
    .Y(_0037_));
 sg13g2_nor2_1 _4608_ (.A(net655),
    .B(net707),
    .Y(_0038_));
 sg13g2_nor2_1 _4609_ (.A(net655),
    .B(net702),
    .Y(_0039_));
 sg13g2_nor2_1 _4610_ (.A(net655),
    .B(net707),
    .Y(_0040_));
 sg13g2_nor2_1 _4611_ (.A(net655),
    .B(net707),
    .Y(_0041_));
 sg13g2_nor2_1 _4612_ (.A(net689),
    .B(net739),
    .Y(_0042_));
 sg13g2_nor2_1 _4613_ (.A(net689),
    .B(net740),
    .Y(_0043_));
 sg13g2_nor2_1 _4614_ (.A(net688),
    .B(net734),
    .Y(_0044_));
 sg13g2_nor2_1 _4615_ (.A(net689),
    .B(net739),
    .Y(_0045_));
 sg13g2_nor2_1 _4616_ (.A(net663),
    .B(net715),
    .Y(_0046_));
 sg13g2_nor2_1 _4617_ (.A(net663),
    .B(net715),
    .Y(_0047_));
 sg13g2_nor2_1 _4618_ (.A(net663),
    .B(net715),
    .Y(_0048_));
 sg13g2_nor2_1 _4619_ (.A(net665),
    .B(net717),
    .Y(_0049_));
 sg13g2_nor2_1 _4620_ (.A(net661),
    .B(net713),
    .Y(_0050_));
 sg13g2_nor2_1 _4621_ (.A(net662),
    .B(net714),
    .Y(_0051_));
 sg13g2_nor2_1 _4622_ (.A(net667),
    .B(net720),
    .Y(_0052_));
 sg13g2_nor2_1 _4623_ (.A(net661),
    .B(net713),
    .Y(_0053_));
 sg13g2_nor2_1 _4624_ (.A(net663),
    .B(net715),
    .Y(_0054_));
 sg13g2_nor2_1 _4625_ (.A(net663),
    .B(net713),
    .Y(_0055_));
 sg13g2_nor2_1 _4626_ (.A(net663),
    .B(net715),
    .Y(_0056_));
 sg13g2_nor2_1 _4627_ (.A(net663),
    .B(net713),
    .Y(_0057_));
 sg13g2_nor2_1 _4628_ (.A(net652),
    .B(net704),
    .Y(_0058_));
 sg13g2_nor2_1 _4629_ (.A(net652),
    .B(net704),
    .Y(_0059_));
 sg13g2_nor2_1 _4630_ (.A(net652),
    .B(net704),
    .Y(_0060_));
 sg13g2_nor2_1 _4631_ (.A(net653),
    .B(net705),
    .Y(_0061_));
 sg13g2_nor2_1 _4632_ (.A(net664),
    .B(net715),
    .Y(_0062_));
 sg13g2_nor2_1 _4633_ (.A(net664),
    .B(net716),
    .Y(_0063_));
 sg13g2_nor2_1 _4634_ (.A(net665),
    .B(net717),
    .Y(_0064_));
 sg13g2_nor2_1 _4635_ (.A(net665),
    .B(net717),
    .Y(_0065_));
 sg13g2_nor2_1 _4636_ (.A(net664),
    .B(net716),
    .Y(_0066_));
 sg13g2_nor2_1 _4637_ (.A(net664),
    .B(net715),
    .Y(_0067_));
 sg13g2_nor2_1 _4638_ (.A(net663),
    .B(net716),
    .Y(_0068_));
 sg13g2_nor2_1 _4639_ (.A(net664),
    .B(net716),
    .Y(_0069_));
 sg13g2_nor2_1 _4640_ (.A(net664),
    .B(net715),
    .Y(_0070_));
 sg13g2_nor2_1 _4641_ (.A(net664),
    .B(net716),
    .Y(_0071_));
 sg13g2_nor2_1 _4642_ (.A(net665),
    .B(net717),
    .Y(_0072_));
 sg13g2_nor2_1 _4643_ (.A(net666),
    .B(net718),
    .Y(_0073_));
 sg13g2_nor2_1 _4644_ (.A(net669),
    .B(net722),
    .Y(_0074_));
 sg13g2_nor2_1 _4645_ (.A(net669),
    .B(net722),
    .Y(_0075_));
 sg13g2_nor2_1 _4646_ (.A(net670),
    .B(net721),
    .Y(_0076_));
 sg13g2_nor2_1 _4647_ (.A(net670),
    .B(net721),
    .Y(_0077_));
 sg13g2_nor2_1 _4648_ (.A(net669),
    .B(net722),
    .Y(_0078_));
 sg13g2_nor2_1 _4649_ (.A(net669),
    .B(net722),
    .Y(_0079_));
 sg13g2_nor2_1 _4650_ (.A(net670),
    .B(net721),
    .Y(_0080_));
 sg13g2_nor2_1 _4651_ (.A(net670),
    .B(net721),
    .Y(_0081_));
 sg13g2_nor2_1 _4652_ (.A(net669),
    .B(net722),
    .Y(_0082_));
 sg13g2_nor2_1 _4653_ (.A(net671),
    .B(net721),
    .Y(_0083_));
 sg13g2_nor2_1 _4654_ (.A(net670),
    .B(net721),
    .Y(_0084_));
 sg13g2_nor2_1 _4655_ (.A(net670),
    .B(net721),
    .Y(_0085_));
 sg13g2_nor2_1 _4656_ (.A(net669),
    .B(net722),
    .Y(_0086_));
 sg13g2_nor2_1 _4657_ (.A(net669),
    .B(net722),
    .Y(_0087_));
 sg13g2_nor2_1 _4658_ (.A(net667),
    .B(net720),
    .Y(_0088_));
 sg13g2_nor2_1 _4659_ (.A(net670),
    .B(net721),
    .Y(_0089_));
 sg13g2_nor2_1 _4660_ (.A(net684),
    .B(net736),
    .Y(_0090_));
 sg13g2_nor2_1 _4661_ (.A(net684),
    .B(net736),
    .Y(_0091_));
 sg13g2_nor2_1 _4662_ (.A(net684),
    .B(net736),
    .Y(_0092_));
 sg13g2_nor2_1 _4663_ (.A(net684),
    .B(net736),
    .Y(_0093_));
 sg13g2_nor2_1 _4664_ (.A(net684),
    .B(net736),
    .Y(_0094_));
 sg13g2_nor2_1 _4665_ (.A(net685),
    .B(net737),
    .Y(_0095_));
 sg13g2_nor2_1 _4666_ (.A(net685),
    .B(net736),
    .Y(_0096_));
 sg13g2_nor2_1 _4667_ (.A(net685),
    .B(net737),
    .Y(_0097_));
 sg13g2_nor2_1 _4668_ (.A(net653),
    .B(net705),
    .Y(_0098_));
 sg13g2_nor2_1 _4669_ (.A(net653),
    .B(net705),
    .Y(_0099_));
 sg13g2_nor2_1 _4670_ (.A(net653),
    .B(net706),
    .Y(_0100_));
 sg13g2_nor2_1 _4671_ (.A(net653),
    .B(net705),
    .Y(_0101_));
 sg13g2_nor2_1 _4672_ (.A(net685),
    .B(net737),
    .Y(_0102_));
 sg13g2_nor2_1 _4673_ (.A(net686),
    .B(net738),
    .Y(_0103_));
 sg13g2_nor2_1 _4674_ (.A(net686),
    .B(net738),
    .Y(_0104_));
 sg13g2_nor2_1 _4675_ (.A(net684),
    .B(net737),
    .Y(_0105_));
 sg13g2_nor2_1 _4676_ (.A(net687),
    .B(net735),
    .Y(_0106_));
 sg13g2_nor2_1 _4677_ (.A(net687),
    .B(net735),
    .Y(_0107_));
 sg13g2_nor2_1 _4678_ (.A(net675),
    .B(net727),
    .Y(_0108_));
 sg13g2_nor2_1 _4679_ (.A(net675),
    .B(net727),
    .Y(_0109_));
 sg13g2_nor2_1 _4680_ (.A(net676),
    .B(net728),
    .Y(_0110_));
 sg13g2_nor2_1 _4681_ (.A(net676),
    .B(net728),
    .Y(_0111_));
 sg13g2_nor2_1 _4682_ (.A(net675),
    .B(net727),
    .Y(_0112_));
 sg13g2_nor2_1 _4683_ (.A(net675),
    .B(net727),
    .Y(_0113_));
 sg13g2_nor2_1 _4684_ (.A(net681),
    .B(net728),
    .Y(_0114_));
 sg13g2_nor2_1 _4685_ (.A(net679),
    .B(net731),
    .Y(_0115_));
 sg13g2_nor2_1 _4686_ (.A(net676),
    .B(net728),
    .Y(_0116_));
 sg13g2_nor2_1 _4687_ (.A(net676),
    .B(net728),
    .Y(_0117_));
 sg13g2_nor2_1 _4688_ (.A(net676),
    .B(net728),
    .Y(_0118_));
 sg13g2_nor2_1 _4689_ (.A(net675),
    .B(net727),
    .Y(_0119_));
 sg13g2_nor2_1 _4690_ (.A(net675),
    .B(net727),
    .Y(_0120_));
 sg13g2_nor2_1 _4691_ (.A(net675),
    .B(net727),
    .Y(_0121_));
 sg13g2_nor2_1 _4692_ (.A(net680),
    .B(net730),
    .Y(_0122_));
 sg13g2_nor2_1 _4693_ (.A(net679),
    .B(net731),
    .Y(_0123_));
 sg13g2_nor2_1 _4694_ (.A(net679),
    .B(net731),
    .Y(_0124_));
 sg13g2_nor2_1 _4695_ (.A(net680),
    .B(net730),
    .Y(_0125_));
 sg13g2_nor2_1 _4696_ (.A(net680),
    .B(net730),
    .Y(_0126_));
 sg13g2_nor2_1 _4697_ (.A(net679),
    .B(net731),
    .Y(_0127_));
 sg13g2_nor2_1 _4698_ (.A(net679),
    .B(net731),
    .Y(_0128_));
 sg13g2_nor2_1 _4699_ (.A(net680),
    .B(net730),
    .Y(_0129_));
 sg13g2_nor2_1 _4700_ (.A(net680),
    .B(net730),
    .Y(_0130_));
 sg13g2_nor2_1 _4701_ (.A(net680),
    .B(net730),
    .Y(_0131_));
 sg13g2_nor2_1 _4702_ (.A(net679),
    .B(net731),
    .Y(_0132_));
 sg13g2_nor2_1 _4703_ (.A(net679),
    .B(net731),
    .Y(_0133_));
 sg13g2_nor2_1 _4704_ (.A(net649),
    .B(net701),
    .Y(_0134_));
 sg13g2_nor2_1 _4705_ (.A(net649),
    .B(net701),
    .Y(_0135_));
 sg13g2_nor2_1 _4706_ (.A(net652),
    .B(net704),
    .Y(_0136_));
 sg13g2_nor2_1 _4707_ (.A(net651),
    .B(net701),
    .Y(_0137_));
 sg13g2_nor2_1 _4708_ (.A(net680),
    .B(net730),
    .Y(_0138_));
 sg13g2_nor2_1 _4709_ (.A(net680),
    .B(net732),
    .Y(_0139_));
 sg13g2_nor2_1 _4710_ (.A(net679),
    .B(net731),
    .Y(_0140_));
 sg13g2_nor2_1 _4711_ (.A(net681),
    .B(net730),
    .Y(_0141_));
 sg13g2_nor2_1 _4712_ (.A(net678),
    .B(net732),
    .Y(_0142_));
 sg13g2_nor2_1 _4713_ (.A(net677),
    .B(net726),
    .Y(_0143_));
 sg13g2_nor2_1 _4714_ (.A(net674),
    .B(net726),
    .Y(_0144_));
 sg13g2_nor2_1 _4715_ (.A(net678),
    .B(net729),
    .Y(_0145_));
 sg13g2_nor2_1 _4716_ (.A(net660),
    .B(net712),
    .Y(_0146_));
 sg13g2_nor2_1 _4717_ (.A(net660),
    .B(net712),
    .Y(_0147_));
 sg13g2_nor2_1 _4718_ (.A(net667),
    .B(net720),
    .Y(_0148_));
 sg13g2_nor2_1 _4719_ (.A(net662),
    .B(net714),
    .Y(_0149_));
 sg13g2_nor2_1 _4720_ (.A(net655),
    .B(net707),
    .Y(_0150_));
 sg13g2_nor2_1 _4721_ (.A(net655),
    .B(net707),
    .Y(_0151_));
 sg13g2_nor2_1 _4722_ (.A(net656),
    .B(net707),
    .Y(_0152_));
 sg13g2_nor2_1 _4723_ (.A(net655),
    .B(net707),
    .Y(_0153_));
 sg13g2_nor2_1 _4724_ (.A(net650),
    .B(net703),
    .Y(_0154_));
 sg13g2_nor2_1 _4725_ (.A(net651),
    .B(net702),
    .Y(_0155_));
 sg13g2_nor2_1 _4726_ (.A(net654),
    .B(net705),
    .Y(_0156_));
 sg13g2_nor2_1 _4727_ (.A(net650),
    .B(net703),
    .Y(_0157_));
 sg13g2_nor2_1 _4728_ (.A(net649),
    .B(net701),
    .Y(_0158_));
 sg13g2_nor2_1 _4729_ (.A(net649),
    .B(net701),
    .Y(_0159_));
 sg13g2_nor2_1 _4730_ (.A(net650),
    .B(net702),
    .Y(_0160_));
 sg13g2_nor2_1 _4731_ (.A(net650),
    .B(net702),
    .Y(_0161_));
 sg13g2_nor2_1 _4732_ (.A(net677),
    .B(net729),
    .Y(_0162_));
 sg13g2_nor2_1 _4733_ (.A(net677),
    .B(net729),
    .Y(_0163_));
 sg13g2_nor2_1 _4734_ (.A(net677),
    .B(net729),
    .Y(_0164_));
 sg13g2_nor2_1 _4735_ (.A(net677),
    .B(net729),
    .Y(_0165_));
 sg13g2_nor2_1 _4736_ (.A(net678),
    .B(net732),
    .Y(_0166_));
 sg13g2_nor2_1 _4737_ (.A(net677),
    .B(net729),
    .Y(_0167_));
 sg13g2_nor2_1 _4738_ (.A(net674),
    .B(net726),
    .Y(_0168_));
 sg13g2_nor2_1 _4739_ (.A(net678),
    .B(net732),
    .Y(_0169_));
 sg13g2_nor2_1 _4740_ (.A(net656),
    .B(net711),
    .Y(_0170_));
 sg13g2_nor2_1 _4741_ (.A(net656),
    .B(net708),
    .Y(_0171_));
 sg13g2_nor2_1 _4742_ (.A(net656),
    .B(net708),
    .Y(_0172_));
 sg13g2_nor2_1 _4743_ (.A(net656),
    .B(net708),
    .Y(_0173_));
 sg13g2_nor2_1 _4744_ (.A(net674),
    .B(net725),
    .Y(_0174_));
 sg13g2_nor2_1 _4745_ (.A(net659),
    .B(net708),
    .Y(_0175_));
 sg13g2_nor2_1 _4746_ (.A(net673),
    .B(net725),
    .Y(_0176_));
 sg13g2_nor2_1 _4747_ (.A(net674),
    .B(net726),
    .Y(_0177_));
 sg13g2_nor2_1 _4748_ (.A(net673),
    .B(net725),
    .Y(_0178_));
 sg13g2_nor2_1 _4749_ (.A(net673),
    .B(net725),
    .Y(_0179_));
 sg13g2_nor2_1 _4750_ (.A(net673),
    .B(net725),
    .Y(_0180_));
 sg13g2_nor2_1 _4751_ (.A(net673),
    .B(net725),
    .Y(_0181_));
 sg13g2_nor2_1 _4752_ (.A(net673),
    .B(net725),
    .Y(_0182_));
 sg13g2_nor2_1 _4753_ (.A(net673),
    .B(net725),
    .Y(_0183_));
 sg13g2_nor2_1 _4754_ (.A(net673),
    .B(net708),
    .Y(_0184_));
 sg13g2_nor2_1 _4755_ (.A(net656),
    .B(net708),
    .Y(_0185_));
 sg13g2_nor2_1 _4756_ (.A(net683),
    .B(net735),
    .Y(_0186_));
 sg13g2_nor2_1 _4757_ (.A(net683),
    .B(net734),
    .Y(_0187_));
 sg13g2_nor2_1 _4758_ (.A(net686),
    .B(net734),
    .Y(_0188_));
 sg13g2_nor2_1 _4759_ (.A(net683),
    .B(net734),
    .Y(_0189_));
 sg13g2_nor2_1 _4760_ (.A(net668),
    .B(net723),
    .Y(_0190_));
 sg13g2_nor2_1 _4761_ (.A(net668),
    .B(net719),
    .Y(_0191_));
 sg13g2_nor2_1 _4762_ (.A(net669),
    .B(net719),
    .Y(_0192_));
 sg13g2_nor2_1 _4763_ (.A(net668),
    .B(net719),
    .Y(_0193_));
 sg13g2_nor2_1 _4764_ (.A(net662),
    .B(net714),
    .Y(_0194_));
 sg13g2_nor2_1 _4765_ (.A(net662),
    .B(net714),
    .Y(_0195_));
 sg13g2_nor2_1 _4766_ (.A(net667),
    .B(net720),
    .Y(_0196_));
 sg13g2_nor2_1 _4767_ (.A(net667),
    .B(net720),
    .Y(_0197_));
 sg13g2_nor2_1 _4768_ (.A(net687),
    .B(net735),
    .Y(_0198_));
 sg13g2_nor2_1 _4769_ (.A(net683),
    .B(net734),
    .Y(_0199_));
 sg13g2_nor2_1 _4770_ (.A(net683),
    .B(net734),
    .Y(_0200_));
 sg13g2_nor2_1 _4771_ (.A(net683),
    .B(net734),
    .Y(_0201_));
 sg13g2_nor2_1 _4772_ (.A(net657),
    .B(net709),
    .Y(_0202_));
 sg13g2_nor2_1 _4773_ (.A(net667),
    .B(net720),
    .Y(_0203_));
 sg13g2_nor2_1 _4774_ (.A(net658),
    .B(net710),
    .Y(_0204_));
 sg13g2_nor2_1 _4775_ (.A(net657),
    .B(net709),
    .Y(_0205_));
 sg13g2_nor2_1 _4776_ (.A(net668),
    .B(net719),
    .Y(_0206_));
 sg13g2_nor2_1 _4777_ (.A(net667),
    .B(net720),
    .Y(_0207_));
 sg13g2_nor2_1 _4778_ (.A(net658),
    .B(net710),
    .Y(_0208_));
 sg13g2_nor2_1 _4779_ (.A(net658),
    .B(net710),
    .Y(_0209_));
 sg13g2_nor2_1 _4780_ (.A(net668),
    .B(net719),
    .Y(_0210_));
 sg13g2_nor2_1 _4781_ (.A(net668),
    .B(net719),
    .Y(_0211_));
 sg13g2_nor2_1 _4782_ (.A(net675),
    .B(net727),
    .Y(_0212_));
 sg13g2_nor2_1 _4783_ (.A(net658),
    .B(net710),
    .Y(_0213_));
 sg13g2_nor2_1 _4784_ (.A(net657),
    .B(net709),
    .Y(_0214_));
 sg13g2_nor2_1 _4785_ (.A(net667),
    .B(net720),
    .Y(_0215_));
 sg13g2_nor2_1 _4786_ (.A(net658),
    .B(net710),
    .Y(_0216_));
 sg13g2_nor2_1 _4787_ (.A(net657),
    .B(net709),
    .Y(_0217_));
 sg13g2_nor2_1 _4788_ (.A(net690),
    .B(net742),
    .Y(_0218_));
 sg13g2_nor2_1 _4789_ (.A(net690),
    .B(net743),
    .Y(_0219_));
 sg13g2_nor2_1 _4790_ (.A(net685),
    .B(net737),
    .Y(_0220_));
 sg13g2_nor2_1 _4791_ (.A(net690),
    .B(net742),
    .Y(_0221_));
 sg13g2_nor2_1 _4792_ (.A(net691),
    .B(net741),
    .Y(_0222_));
 sg13g2_nor2_1 _4793_ (.A(net690),
    .B(net741),
    .Y(_0223_));
 sg13g2_nor2_1 _4794_ (.A(net691),
    .B(net741),
    .Y(_0224_));
 sg13g2_nor2_1 _4795_ (.A(net690),
    .B(net742),
    .Y(_0225_));
 sg13g2_nor2_1 _4796_ (.A(net690),
    .B(net742),
    .Y(_0226_));
 sg13g2_nor2_1 _4797_ (.A(net692),
    .B(net742),
    .Y(_0227_));
 sg13g2_nor2_1 _4798_ (.A(net691),
    .B(net742),
    .Y(_0228_));
 sg13g2_nor2_1 _4799_ (.A(net691),
    .B(net742),
    .Y(_0229_));
 sg13g2_nor2_1 _4800_ (.A(net690),
    .B(net741),
    .Y(_0230_));
 sg13g2_nor2_1 _4801_ (.A(net691),
    .B(net741),
    .Y(_0231_));
 sg13g2_nor2_1 _4802_ (.A(net691),
    .B(net741),
    .Y(_0232_));
 sg13g2_nor2_1 _4803_ (.A(net690),
    .B(net741),
    .Y(_0233_));
 sg13g2_nor2_1 _4804_ (.A(net660),
    .B(net712),
    .Y(_0234_));
 sg13g2_nor2_1 _4805_ (.A(net660),
    .B(net712),
    .Y(_0235_));
 sg13g2_nor2_1 _4806_ (.A(net653),
    .B(net705),
    .Y(_0236_));
 sg13g2_nor2_1 _4807_ (.A(net660),
    .B(net712),
    .Y(_0237_));
 sg13g2_nor2_1 _4808_ (.A(net688),
    .B(net740),
    .Y(_0238_));
 sg13g2_nor2_1 _4809_ (.A(net689),
    .B(net739),
    .Y(_0239_));
 sg13g2_nor2_1 _4810_ (.A(net688),
    .B(net740),
    .Y(_0240_));
 sg13g2_nor2_1 _4811_ (.A(net689),
    .B(net739),
    .Y(_0241_));
 sg13g2_nor2_1 _4812_ (.A(net689),
    .B(net739),
    .Y(_0242_));
 sg13g2_nor2_1 _4813_ (.A(net689),
    .B(net743),
    .Y(_0243_));
 sg13g2_nor2_1 _4814_ (.A(net688),
    .B(net740),
    .Y(_0244_));
 sg13g2_nor2_1 _4815_ (.A(net688),
    .B(net740),
    .Y(_0245_));
 sg13g2_nor2_1 _4816_ (.A(net688),
    .B(net740),
    .Y(_0246_));
 sg13g2_nor2_1 _4817_ (.A(net691),
    .B(net741),
    .Y(_0247_));
 sg13g2_nor2_1 _4818_ (.A(net688),
    .B(net735),
    .Y(_0248_));
 sg13g2_nor2_1 _4819_ (.A(net688),
    .B(net740),
    .Y(_0249_));
 sg13g2_nor2_1 _4820_ (.A(net652),
    .B(net704),
    .Y(_0250_));
 sg13g2_nor2_1 _4821_ (.A(net653),
    .B(net705),
    .Y(_0251_));
 sg13g2_nor2_1 _4822_ (.A(net654),
    .B(net706),
    .Y(_0252_));
 sg13g2_nor2_1 _4823_ (.A(net652),
    .B(net704),
    .Y(_0253_));
 sg13g2_nor2_1 _4824_ (.A(net655),
    .B(net707),
    .Y(_0254_));
 sg13g2_nor2_1 _4825_ (.A(net656),
    .B(net708),
    .Y(_0255_));
 sg13g2_nor2_1 _4826_ (.A(net657),
    .B(net709),
    .Y(_0256_));
 sg13g2_nor2_1 _4827_ (.A(net657),
    .B(net709),
    .Y(_0257_));
 sg13g2_nor2_1 _4828_ (.A(_2064_),
    .B(_2068_),
    .Y(_0613_));
 sg13g2_nor2_1 _4829_ (.A(_2064_),
    .B(_2068_),
    .Y(_0614_));
 sg13g2_nor2_1 _4830_ (.A(net650),
    .B(net702),
    .Y(_0258_));
 sg13g2_nor2_1 _4831_ (.A(net650),
    .B(net702),
    .Y(_0259_));
 sg13g2_nor2_1 _4832_ (.A(net650),
    .B(net702),
    .Y(_0260_));
 sg13g2_nor2_1 _4833_ (.A(net650),
    .B(net702),
    .Y(_0261_));
 sg13g2_dfrbpq_1 _4834_ (.RESET_B(net261),
    .D(_0263_),
    .Q(\tmds_green.dc_balancing_reg[0] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4835_ (.RESET_B(net158),
    .D(_0264_),
    .Q(\tmds_blue.dc_balancing_reg[0] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _4836_ (.RESET_B(net156),
    .D(_0265_),
    .Q(\clockdiv.q1 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _4837_ (.RESET_B(net155),
    .D(_0266_),
    .Q(\clockdiv.q2 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _4838_ (.RESET_B(net154),
    .D(net743),
    .Q(\clockdiv.q2temp ),
    .CLK(net405));
 sg13g2_dfrbpq_1 _4839_ (.RESET_B(net153),
    .D(_0267_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][0] ),
    .CLK(_0006_));
 sg13g2_dfrbpq_1 _4840_ (.RESET_B(net151),
    .D(_0268_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][1] ),
    .CLK(_0007_));
 sg13g2_dfrbpq_1 _4841_ (.RESET_B(net149),
    .D(_0269_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][2] ),
    .CLK(_0008_));
 sg13g2_dfrbpq_1 _4842_ (.RESET_B(net147),
    .D(_0270_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[39][3] ),
    .CLK(_0009_));
 sg13g2_dfrbpq_1 _4843_ (.RESET_B(net145),
    .D(_0271_),
    .Q(\green_tmds_par[0] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _4844_ (.RESET_B(net144),
    .D(_0272_),
    .Q(\green_tmds_par[1] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _4845_ (.RESET_B(net143),
    .D(_0273_),
    .Q(\green_tmds_par[7] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _4846_ (.RESET_B(net142),
    .D(_0274_),
    .Q(\red_tmds_par[0] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4847_ (.RESET_B(net141),
    .D(_0275_),
    .Q(\red_tmds_par[1] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _4848_ (.RESET_B(net140),
    .D(_0276_),
    .Q(\red_tmds_par[3] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4849_ (.RESET_B(net139),
    .D(_0277_),
    .Q(\red_tmds_par[5] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4850_ (.RESET_B(net138),
    .D(_0278_),
    .Q(\red_tmds_par[7] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4851_ (.RESET_B(net137),
    .D(_0279_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][0] ),
    .CLK(_0010_));
 sg13g2_dfrbpq_1 _4852_ (.RESET_B(net135),
    .D(_0280_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][1] ),
    .CLK(_0011_));
 sg13g2_dfrbpq_1 _4853_ (.RESET_B(net133),
    .D(_0281_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][2] ),
    .CLK(_0012_));
 sg13g2_dfrbpq_1 _4854_ (.RESET_B(net131),
    .D(_0282_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[59][3] ),
    .CLK(_0013_));
 sg13g2_dfrbpq_1 _4855_ (.RESET_B(net129),
    .D(_0283_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][0] ),
    .CLK(_0014_));
 sg13g2_dfrbpq_1 _4856_ (.RESET_B(net127),
    .D(_0284_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][1] ),
    .CLK(_0015_));
 sg13g2_dfrbpq_1 _4857_ (.RESET_B(net125),
    .D(_0285_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][2] ),
    .CLK(_0016_));
 sg13g2_dfrbpq_1 _4858_ (.RESET_B(net123),
    .D(_0286_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[6][3] ),
    .CLK(_0017_));
 sg13g2_dfrbpq_1 _4859_ (.RESET_B(net121),
    .D(_0287_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][0] ),
    .CLK(_0018_));
 sg13g2_dfrbpq_1 _4860_ (.RESET_B(net119),
    .D(_0288_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][1] ),
    .CLK(_0019_));
 sg13g2_dfrbpq_1 _4861_ (.RESET_B(net117),
    .D(_0289_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][2] ),
    .CLK(_0020_));
 sg13g2_dfrbpq_1 _4862_ (.RESET_B(net115),
    .D(_0290_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[49][3] ),
    .CLK(_0021_));
 sg13g2_dfrbpq_1 _4863_ (.RESET_B(net113),
    .D(_0291_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][0] ),
    .CLK(_0022_));
 sg13g2_dfrbpq_1 _4864_ (.RESET_B(net111),
    .D(_0292_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][1] ),
    .CLK(_0023_));
 sg13g2_dfrbpq_1 _4865_ (.RESET_B(net109),
    .D(_0293_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][2] ),
    .CLK(_0024_));
 sg13g2_dfrbpq_1 _4866_ (.RESET_B(net107),
    .D(_0294_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[9][3] ),
    .CLK(_0025_));
 sg13g2_dfrbpq_1 _4867_ (.RESET_B(net105),
    .D(_0295_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][0] ),
    .CLK(_0026_));
 sg13g2_dfrbpq_1 _4868_ (.RESET_B(net103),
    .D(_0296_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][1] ),
    .CLK(_0027_));
 sg13g2_dfrbpq_1 _4869_ (.RESET_B(net101),
    .D(_0297_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][2] ),
    .CLK(_0028_));
 sg13g2_dfrbpq_1 _4870_ (.RESET_B(net99),
    .D(_0298_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[63][3] ),
    .CLK(_0029_));
 sg13g2_dfrbpq_2 _4871_ (.RESET_B(net97),
    .D(_0299_),
    .Q(\videogen.fancy_shader.video_x[0] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4872_ (.RESET_B(net96),
    .D(_0300_),
    .Q(\videogen.fancy_shader.video_x[1] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4873_ (.RESET_B(net95),
    .D(_0301_),
    .Q(\videogen.fancy_shader.video_x[2] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4874_ (.RESET_B(net94),
    .D(_0302_),
    .Q(\videogen.fancy_shader.video_x[3] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4875_ (.RESET_B(net93),
    .D(_0303_),
    .Q(\videogen.fancy_shader.video_x[4] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4876_ (.RESET_B(net92),
    .D(_0304_),
    .Q(\videogen.fancy_shader.video_x[5] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4877_ (.RESET_B(net91),
    .D(_0305_),
    .Q(\videogen.fancy_shader.video_x[6] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4878_ (.RESET_B(net90),
    .D(_0306_),
    .Q(\videogen.fancy_shader.video_x[7] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4879_ (.RESET_B(net89),
    .D(_0307_),
    .Q(\videogen.fancy_shader.video_x[8] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4880_ (.RESET_B(net88),
    .D(_0308_),
    .Q(\videogen.fancy_shader.video_x[9] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4881_ (.RESET_B(net87),
    .D(_0309_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][0] ),
    .CLK(_0030_));
 sg13g2_dfrbpq_1 _4882_ (.RESET_B(net85),
    .D(_0310_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][1] ),
    .CLK(_0031_));
 sg13g2_dfrbpq_1 _4883_ (.RESET_B(net83),
    .D(_0311_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][2] ),
    .CLK(_0032_));
 sg13g2_dfrbpq_1 _4884_ (.RESET_B(net81),
    .D(_0312_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[0][3] ),
    .CLK(_0033_));
 sg13g2_dfrbpq_1 _4885_ (.RESET_B(net79),
    .D(_0313_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][0] ),
    .CLK(_0034_));
 sg13g2_dfrbpq_1 _4886_ (.RESET_B(net77),
    .D(_0314_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][1] ),
    .CLK(_0035_));
 sg13g2_dfrbpq_1 _4887_ (.RESET_B(net75),
    .D(_0315_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][2] ),
    .CLK(_0036_));
 sg13g2_dfrbpq_1 _4888_ (.RESET_B(net73),
    .D(_0316_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[29][3] ),
    .CLK(_0037_));
 sg13g2_dfrbpq_1 _4889_ (.RESET_B(net71),
    .D(_0317_),
    .Q(\tmds_blue.vsync ),
    .CLK(net636));
 sg13g2_dfrbpq_1 _4890_ (.RESET_B(net70),
    .D(_0318_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[0] ),
    .CLK(net631));
 sg13g2_dfrbpq_1 _4891_ (.RESET_B(net68),
    .D(_0319_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[1] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4892_ (.RESET_B(net66),
    .D(_0320_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[2] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4893_ (.RESET_B(net64),
    .D(_0321_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[3] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4894_ (.RESET_B(net62),
    .D(_0322_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[4] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4895_ (.RESET_B(net60),
    .D(_0323_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_pix[5] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4896_ (.RESET_B(net58),
    .D(_0324_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ),
    .CLK(net630));
 sg13g2_dfrbpq_2 _4897_ (.RESET_B(net56),
    .D(_0325_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[1] ),
    .CLK(net631));
 sg13g2_dfrbpq_2 _4898_ (.RESET_B(net54),
    .D(_0326_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .CLK(net630));
 sg13g2_dfrbpq_2 _4899_ (.RESET_B(net52),
    .D(_0327_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .CLK(net630));
 sg13g2_dfrbpq_2 _4900_ (.RESET_B(net50),
    .D(_0328_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .CLK(net630));
 sg13g2_dfrbpq_2 _4901_ (.RESET_B(net48),
    .D(_0329_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .CLK(net648));
 sg13g2_dfrbpq_1 _4902_ (.RESET_B(net46),
    .D(_0330_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[0] ),
    .CLK(net630));
 sg13g2_dfrbpq_1 _4903_ (.RESET_B(net44),
    .D(_0331_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[1] ),
    .CLK(net630));
 sg13g2_dfrbpq_1 _4904_ (.RESET_B(net42),
    .D(_0332_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[2] ),
    .CLK(net630));
 sg13g2_dfrbpq_1 _4905_ (.RESET_B(net40),
    .D(_0333_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.v_counter[3] ),
    .CLK(net630));
 sg13g2_dfrbpq_1 _4906_ (.RESET_B(net38),
    .D(_0334_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[0] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _4907_ (.RESET_B(net36),
    .D(_0335_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[1] ),
    .CLK(net635));
 sg13g2_dfrbpq_2 _4908_ (.RESET_B(net34),
    .D(_0336_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[2] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _4909_ (.RESET_B(net32),
    .D(_0337_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.h_counter[3] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _4910_ (.RESET_B(net404),
    .D(_0338_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][0] ),
    .CLK(_0038_));
 sg13g2_dfrbpq_1 _4911_ (.RESET_B(net400),
    .D(_0339_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][1] ),
    .CLK(_0039_));
 sg13g2_dfrbpq_1 _4912_ (.RESET_B(net398),
    .D(_0340_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][2] ),
    .CLK(_0040_));
 sg13g2_dfrbpq_1 _4913_ (.RESET_B(net396),
    .D(_0341_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[12][3] ),
    .CLK(_0041_));
 sg13g2_dfrbpq_1 _4914_ (.RESET_B(net394),
    .D(_0342_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][0] ),
    .CLK(_0042_));
 sg13g2_dfrbpq_1 _4915_ (.RESET_B(net392),
    .D(_0343_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][1] ),
    .CLK(_0043_));
 sg13g2_dfrbpq_1 _4916_ (.RESET_B(net390),
    .D(_0344_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][2] ),
    .CLK(_0044_));
 sg13g2_dfrbpq_1 _4917_ (.RESET_B(net388),
    .D(_0345_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[19][3] ),
    .CLK(_0045_));
 sg13g2_dfrbpq_2 _4918_ (.RESET_B(net386),
    .D(_0346_),
    .Q(\videogen.fancy_shader.n646[0] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4919_ (.RESET_B(net384),
    .D(_0347_),
    .Q(\videogen.fancy_shader.n646[1] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4920_ (.RESET_B(net382),
    .D(_0348_),
    .Q(\videogen.fancy_shader.n646[2] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4921_ (.RESET_B(net380),
    .D(_0349_),
    .Q(\videogen.fancy_shader.n646[3] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4922_ (.RESET_B(net378),
    .D(_0350_),
    .Q(\videogen.fancy_shader.n646[4] ),
    .CLK(net647));
 sg13g2_dfrbpq_2 _4923_ (.RESET_B(net376),
    .D(_0351_),
    .Q(\videogen.fancy_shader.n646[5] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4924_ (.RESET_B(net374),
    .D(_0352_),
    .Q(\videogen.fancy_shader.n646[6] ),
    .CLK(net634));
 sg13g2_dfrbpq_2 _4925_ (.RESET_B(net372),
    .D(_0353_),
    .Q(\videogen.fancy_shader.n646[7] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4926_ (.RESET_B(net370),
    .D(_0354_),
    .Q(\videogen.fancy_shader.n646[8] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4927_ (.RESET_B(net368),
    .D(_0355_),
    .Q(\videogen.fancy_shader.n646[9] ),
    .CLK(net634));
 sg13g2_dfrbpq_1 _4928_ (.RESET_B(net366),
    .D(_0356_),
    .Q(\videogen.fancy_shader.video_y[0] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4929_ (.RESET_B(net364),
    .D(_0357_),
    .Q(\videogen.fancy_shader.video_y[1] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4930_ (.RESET_B(net362),
    .D(_0358_),
    .Q(\videogen.fancy_shader.video_y[2] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4931_ (.RESET_B(net360),
    .D(_0359_),
    .Q(\videogen.fancy_shader.video_y[3] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4932_ (.RESET_B(net358),
    .D(_0360_),
    .Q(\videogen.fancy_shader.video_y[4] ),
    .CLK(net633));
 sg13g2_dfrbpq_2 _4933_ (.RESET_B(net356),
    .D(_0361_),
    .Q(\videogen.fancy_shader.video_y[5] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4934_ (.RESET_B(net354),
    .D(_0362_),
    .Q(\videogen.fancy_shader.video_y[6] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4935_ (.RESET_B(net352),
    .D(_0363_),
    .Q(\videogen.fancy_shader.video_y[7] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4936_ (.RESET_B(net350),
    .D(_0364_),
    .Q(\videogen.fancy_shader.video_y[8] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4937_ (.RESET_B(net348),
    .D(_0365_),
    .Q(\videogen.fancy_shader.video_y[9] ),
    .CLK(net632));
 sg13g2_dfrbpq_2 _4938_ (.RESET_B(net346),
    .D(_0366_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[0] ),
    .CLK(net639));
 sg13g2_dfrbpq_2 _4939_ (.RESET_B(net345),
    .D(_0367_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[1] ),
    .CLK(net639));
 sg13g2_dfrbpq_1 _4940_ (.RESET_B(net344),
    .D(_0368_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[2] ),
    .CLK(net639));
 sg13g2_dfrbpq_1 _4941_ (.RESET_B(net343),
    .D(_0369_),
    .Q(\videogen.test_lut_thingy.gol_counter_reg[3] ),
    .CLK(net639));
 sg13g2_dfrbpq_2 _4942_ (.RESET_B(net342),
    .D(_0370_),
    .Q(hsync),
    .CLK(net639));
 sg13g2_dfrbpq_1 _4943_ (.RESET_B(net341),
    .D(_0371_),
    .Q(display_enable),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4944_ (.RESET_B(net340),
    .D(_0372_),
    .Q(\tmds_blue.n193 ),
    .CLK(net636));
 sg13g2_dfrbpq_1 _4945_ (.RESET_B(net339),
    .D(_0373_),
    .Q(\tmds_blue.n100 ),
    .CLK(net636));
 sg13g2_dfrbpq_1 _4946_ (.RESET_B(net338),
    .D(_0374_),
    .Q(\tmds_blue.n126 ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4947_ (.RESET_B(net337),
    .D(_0375_),
    .Q(\tmds_blue.n132 ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4948_ (.RESET_B(net336),
    .D(_0376_),
    .Q(\tmds_green.n100 ),
    .CLK(net636));
 sg13g2_dfrbpq_2 _4949_ (.RESET_B(net335),
    .D(_0377_),
    .Q(\tmds_green.n126 ),
    .CLK(net643));
 sg13g2_dfrbpq_2 _4950_ (.RESET_B(net334),
    .D(_0378_),
    .Q(\tmds_green.n132 ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _4951_ (.RESET_B(net333),
    .D(_0379_),
    .Q(\tmds_red.n102 ),
    .CLK(net641));
 sg13g2_dfrbpq_2 _4952_ (.RESET_B(net332),
    .D(_0380_),
    .Q(\tmds_red.n100 ),
    .CLK(net642));
 sg13g2_dfrbpq_2 _4953_ (.RESET_B(net331),
    .D(_0381_),
    .Q(\tmds_red.n114 ),
    .CLK(net642));
 sg13g2_dfrbpq_2 _4954_ (.RESET_B(net330),
    .D(_0382_),
    .Q(\tmds_red.n126 ),
    .CLK(net642));
 sg13g2_dfrbpq_2 _4955_ (.RESET_B(net329),
    .D(_0383_),
    .Q(\tmds_red.n132 ),
    .CLK(net642));
 sg13g2_dfrbpq_1 _4956_ (.RESET_B(net328),
    .D(_0384_),
    .Q(\red_tmds_par[2] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4957_ (.RESET_B(net327),
    .D(_0385_),
    .Q(\red_tmds_par[4] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4958_ (.RESET_B(net326),
    .D(_0386_),
    .Q(\red_tmds_par[6] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4959_ (.RESET_B(net325),
    .D(_0387_),
    .Q(\red_tmds_par[8] ),
    .CLK(net636));
 sg13g2_dfrbpq_1 _4960_ (.RESET_B(net324),
    .D(_0388_),
    .Q(\red_tmds_par[9] ),
    .CLK(net641));
 sg13g2_dfrbpq_1 _4961_ (.RESET_B(net323),
    .D(_0389_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][0] ),
    .CLK(_0046_));
 sg13g2_dfrbpq_1 _4962_ (.RESET_B(net321),
    .D(_0390_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][1] ),
    .CLK(_0047_));
 sg13g2_dfrbpq_1 _4963_ (.RESET_B(net319),
    .D(_0391_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][2] ),
    .CLK(_0048_));
 sg13g2_dfrbpq_1 _4964_ (.RESET_B(net317),
    .D(_0392_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[62][3] ),
    .CLK(_0049_));
 sg13g2_dfrbpq_1 _4965_ (.RESET_B(net315),
    .D(_0393_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][0] ),
    .CLK(_0050_));
 sg13g2_dfrbpq_1 _4966_ (.RESET_B(net313),
    .D(_0394_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][1] ),
    .CLK(_0051_));
 sg13g2_dfrbpq_1 _4967_ (.RESET_B(net311),
    .D(_0395_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][2] ),
    .CLK(_0052_));
 sg13g2_dfrbpq_1 _4968_ (.RESET_B(net309),
    .D(_0396_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[61][3] ),
    .CLK(_0053_));
 sg13g2_dfrbpq_1 _4969_ (.RESET_B(net307),
    .D(_0397_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][0] ),
    .CLK(_0054_));
 sg13g2_dfrbpq_1 _4970_ (.RESET_B(net305),
    .D(_0398_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][1] ),
    .CLK(_0055_));
 sg13g2_dfrbpq_1 _4971_ (.RESET_B(net303),
    .D(_0399_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][2] ),
    .CLK(_0056_));
 sg13g2_dfrbpq_1 _4972_ (.RESET_B(net301),
    .D(_0400_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[60][3] ),
    .CLK(_0057_));
 sg13g2_dfrbpq_1 _4973_ (.RESET_B(net300),
    .D(_0401_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][0] ),
    .CLK(_0058_));
 sg13g2_dfrbpq_1 _4974_ (.RESET_B(net298),
    .D(_0402_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][1] ),
    .CLK(_0059_));
 sg13g2_dfrbpq_1 _4975_ (.RESET_B(net296),
    .D(_0403_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][2] ),
    .CLK(_0060_));
 sg13g2_dfrbpq_1 _4976_ (.RESET_B(net294),
    .D(_0404_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[5][3] ),
    .CLK(_0061_));
 sg13g2_dfrbpq_1 _4977_ (.RESET_B(net292),
    .D(_0405_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][0] ),
    .CLK(_0062_));
 sg13g2_dfrbpq_1 _4978_ (.RESET_B(net290),
    .D(_0406_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][1] ),
    .CLK(_0063_));
 sg13g2_dfrbpq_1 _4979_ (.RESET_B(net288),
    .D(_0407_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][2] ),
    .CLK(_0064_));
 sg13g2_dfrbpq_1 _4980_ (.RESET_B(net286),
    .D(_0408_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[58][3] ),
    .CLK(_0065_));
 sg13g2_dfrbpq_1 _4981_ (.RESET_B(net284),
    .D(_0409_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][0] ),
    .CLK(_0066_));
 sg13g2_dfrbpq_1 _4982_ (.RESET_B(net282),
    .D(_0410_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][1] ),
    .CLK(_0067_));
 sg13g2_dfrbpq_1 _4983_ (.RESET_B(net280),
    .D(_0411_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][2] ),
    .CLK(_0068_));
 sg13g2_dfrbpq_1 _4984_ (.RESET_B(net278),
    .D(_0412_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[57][3] ),
    .CLK(_0069_));
 sg13g2_dfrbpq_1 _4985_ (.RESET_B(net276),
    .D(_0413_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][0] ),
    .CLK(_0070_));
 sg13g2_dfrbpq_1 _4986_ (.RESET_B(net274),
    .D(_0414_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][1] ),
    .CLK(_0071_));
 sg13g2_dfrbpq_1 _4987_ (.RESET_B(net272),
    .D(_0415_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][2] ),
    .CLK(_0072_));
 sg13g2_dfrbpq_1 _4988_ (.RESET_B(net270),
    .D(_0416_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[56][3] ),
    .CLK(_0073_));
 sg13g2_dfrbpq_1 _4989_ (.RESET_B(net269),
    .D(_0417_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][0] ),
    .CLK(_0074_));
 sg13g2_dfrbpq_1 _4990_ (.RESET_B(net267),
    .D(_0418_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][1] ),
    .CLK(_0075_));
 sg13g2_dfrbpq_1 _4991_ (.RESET_B(net265),
    .D(_0419_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][2] ),
    .CLK(_0076_));
 sg13g2_dfrbpq_1 _4992_ (.RESET_B(net259),
    .D(_0420_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[55][3] ),
    .CLK(_0077_));
 sg13g2_dfrbpq_1 _4993_ (.RESET_B(net257),
    .D(_0421_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][0] ),
    .CLK(_0078_));
 sg13g2_dfrbpq_1 _4994_ (.RESET_B(net255),
    .D(_0422_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][1] ),
    .CLK(_0079_));
 sg13g2_dfrbpq_1 _4995_ (.RESET_B(net253),
    .D(_0423_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][2] ),
    .CLK(_0080_));
 sg13g2_dfrbpq_1 _4996_ (.RESET_B(net251),
    .D(_0424_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[54][3] ),
    .CLK(_0081_));
 sg13g2_dfrbpq_1 _4997_ (.RESET_B(net249),
    .D(_0425_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][0] ),
    .CLK(_0082_));
 sg13g2_dfrbpq_1 _4998_ (.RESET_B(net247),
    .D(_0426_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][1] ),
    .CLK(_0083_));
 sg13g2_dfrbpq_1 _4999_ (.RESET_B(net245),
    .D(_0427_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][2] ),
    .CLK(_0084_));
 sg13g2_dfrbpq_1 _5000_ (.RESET_B(net243),
    .D(_0428_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[53][3] ),
    .CLK(_0085_));
 sg13g2_dfrbpq_1 _5001_ (.RESET_B(net241),
    .D(_0429_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][0] ),
    .CLK(_0086_));
 sg13g2_dfrbpq_1 _5002_ (.RESET_B(net239),
    .D(_0430_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][1] ),
    .CLK(_0087_));
 sg13g2_dfrbpq_1 _5003_ (.RESET_B(net237),
    .D(_0431_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][2] ),
    .CLK(_0088_));
 sg13g2_dfrbpq_1 _5004_ (.RESET_B(net235),
    .D(_0432_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[52][3] ),
    .CLK(_0089_));
 sg13g2_dfrbpq_1 _5005_ (.RESET_B(net234),
    .D(_0433_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][0] ),
    .CLK(_0090_));
 sg13g2_dfrbpq_1 _5006_ (.RESET_B(net232),
    .D(_0434_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][1] ),
    .CLK(_0091_));
 sg13g2_dfrbpq_1 _5007_ (.RESET_B(net230),
    .D(_0435_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][2] ),
    .CLK(_0092_));
 sg13g2_dfrbpq_1 _5008_ (.RESET_B(net228),
    .D(_0436_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[51][3] ),
    .CLK(_0093_));
 sg13g2_dfrbpq_1 _5009_ (.RESET_B(net226),
    .D(_0437_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][0] ),
    .CLK(_0094_));
 sg13g2_dfrbpq_1 _5010_ (.RESET_B(net224),
    .D(_0438_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][1] ),
    .CLK(_0095_));
 sg13g2_dfrbpq_1 _5011_ (.RESET_B(net222),
    .D(_0439_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][2] ),
    .CLK(_0096_));
 sg13g2_dfrbpq_1 _5012_ (.RESET_B(net220),
    .D(_0440_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[50][3] ),
    .CLK(_0097_));
 sg13g2_dfrbpq_1 _5013_ (.RESET_B(net218),
    .D(_0441_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][0] ),
    .CLK(_0098_));
 sg13g2_dfrbpq_1 _5014_ (.RESET_B(net216),
    .D(_0442_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][1] ),
    .CLK(_0099_));
 sg13g2_dfrbpq_1 _5015_ (.RESET_B(net214),
    .D(_0443_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][2] ),
    .CLK(_0100_));
 sg13g2_dfrbpq_1 _5016_ (.RESET_B(net212),
    .D(_0444_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[4][3] ),
    .CLK(_0101_));
 sg13g2_dfrbpq_1 _5017_ (.RESET_B(net210),
    .D(_0445_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][0] ),
    .CLK(_0102_));
 sg13g2_dfrbpq_1 _5018_ (.RESET_B(net208),
    .D(_0446_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][1] ),
    .CLK(_0103_));
 sg13g2_dfrbpq_1 _5019_ (.RESET_B(net206),
    .D(_0447_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][2] ),
    .CLK(_0104_));
 sg13g2_dfrbpq_1 _5020_ (.RESET_B(net204),
    .D(_0448_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[48][3] ),
    .CLK(_0105_));
 sg13g2_dfrbpq_1 _5021_ (.RESET_B(net202),
    .D(_0449_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][0] ),
    .CLK(_0106_));
 sg13g2_dfrbpq_1 _5022_ (.RESET_B(net200),
    .D(_0450_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][1] ),
    .CLK(_0107_));
 sg13g2_dfrbpq_1 _5023_ (.RESET_B(net198),
    .D(_0451_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][2] ),
    .CLK(_0108_));
 sg13g2_dfrbpq_1 _5024_ (.RESET_B(net196),
    .D(_0452_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[47][3] ),
    .CLK(_0109_));
 sg13g2_dfrbpq_1 _5025_ (.RESET_B(net194),
    .D(_0453_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][0] ),
    .CLK(_0110_));
 sg13g2_dfrbpq_1 _5026_ (.RESET_B(net192),
    .D(_0454_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][1] ),
    .CLK(_0111_));
 sg13g2_dfrbpq_1 _5027_ (.RESET_B(net190),
    .D(_0455_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][2] ),
    .CLK(_0112_));
 sg13g2_dfrbpq_1 _5028_ (.RESET_B(net188),
    .D(_0456_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[46][3] ),
    .CLK(_0113_));
 sg13g2_dfrbpq_1 _5029_ (.RESET_B(net186),
    .D(_0457_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][0] ),
    .CLK(_0114_));
 sg13g2_dfrbpq_1 _5030_ (.RESET_B(net184),
    .D(_0458_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][1] ),
    .CLK(_0115_));
 sg13g2_dfrbpq_1 _5031_ (.RESET_B(net182),
    .D(_0459_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][2] ),
    .CLK(_0116_));
 sg13g2_dfrbpq_1 _5032_ (.RESET_B(net180),
    .D(_0460_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[45][3] ),
    .CLK(_0117_));
 sg13g2_dfrbpq_1 _5033_ (.RESET_B(net178),
    .D(_0461_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][0] ),
    .CLK(_0118_));
 sg13g2_dfrbpq_1 _5034_ (.RESET_B(net176),
    .D(_0462_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][1] ),
    .CLK(_0119_));
 sg13g2_dfrbpq_1 _5035_ (.RESET_B(net174),
    .D(_0463_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][2] ),
    .CLK(_0120_));
 sg13g2_dfrbpq_1 _5036_ (.RESET_B(net172),
    .D(_0464_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[44][3] ),
    .CLK(_0121_));
 sg13g2_dfrbpq_1 _5037_ (.RESET_B(net170),
    .D(_0465_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][0] ),
    .CLK(_0122_));
 sg13g2_dfrbpq_1 _5038_ (.RESET_B(net168),
    .D(_0466_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][1] ),
    .CLK(_0123_));
 sg13g2_dfrbpq_1 _5039_ (.RESET_B(net166),
    .D(_0467_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][2] ),
    .CLK(_0124_));
 sg13g2_dfrbpq_1 _5040_ (.RESET_B(net164),
    .D(_0468_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[43][3] ),
    .CLK(_0125_));
 sg13g2_dfrbpq_1 _5041_ (.RESET_B(net162),
    .D(_0469_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][0] ),
    .CLK(_0126_));
 sg13g2_dfrbpq_1 _5042_ (.RESET_B(net160),
    .D(_0470_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][1] ),
    .CLK(_0127_));
 sg13g2_dfrbpq_1 _5043_ (.RESET_B(net157),
    .D(_0471_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][2] ),
    .CLK(_0128_));
 sg13g2_dfrbpq_1 _5044_ (.RESET_B(net150),
    .D(_0472_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[42][3] ),
    .CLK(_0129_));
 sg13g2_dfrbpq_1 _5045_ (.RESET_B(net146),
    .D(_0473_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][0] ),
    .CLK(_0130_));
 sg13g2_dfrbpq_1 _5046_ (.RESET_B(net134),
    .D(_0474_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][1] ),
    .CLK(_0131_));
 sg13g2_dfrbpq_1 _5047_ (.RESET_B(net130),
    .D(_0475_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][2] ),
    .CLK(_0132_));
 sg13g2_dfrbpq_1 _5048_ (.RESET_B(net126),
    .D(_0476_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[41][3] ),
    .CLK(_0133_));
 sg13g2_dfrbpq_1 _5049_ (.RESET_B(net122),
    .D(_0477_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][0] ),
    .CLK(_0134_));
 sg13g2_dfrbpq_1 _5050_ (.RESET_B(net118),
    .D(_0478_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][1] ),
    .CLK(_0135_));
 sg13g2_dfrbpq_1 _5051_ (.RESET_B(net114),
    .D(_0479_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][2] ),
    .CLK(_0136_));
 sg13g2_dfrbpq_1 _5052_ (.RESET_B(net110),
    .D(_0480_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[8][3] ),
    .CLK(_0137_));
 sg13g2_dfrbpq_1 _5053_ (.RESET_B(net106),
    .D(_0481_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][0] ),
    .CLK(_0138_));
 sg13g2_dfrbpq_1 _5054_ (.RESET_B(net102),
    .D(_0482_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][1] ),
    .CLK(_0139_));
 sg13g2_dfrbpq_1 _5055_ (.RESET_B(net98),
    .D(_0483_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][2] ),
    .CLK(_0140_));
 sg13g2_dfrbpq_1 _5056_ (.RESET_B(net84),
    .D(_0484_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[40][3] ),
    .CLK(_0141_));
 sg13g2_dfrbpq_1 _5057_ (.RESET_B(net80),
    .D(_0485_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][0] ),
    .CLK(_0142_));
 sg13g2_dfrbpq_1 _5058_ (.RESET_B(net76),
    .D(_0486_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][1] ),
    .CLK(_0143_));
 sg13g2_dfrbpq_1 _5059_ (.RESET_B(net72),
    .D(_0487_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][2] ),
    .CLK(_0144_));
 sg13g2_dfrbpq_1 _5060_ (.RESET_B(net67),
    .D(_0488_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[38][3] ),
    .CLK(_0145_));
 sg13g2_dfrbpq_1 _5061_ (.RESET_B(net63),
    .D(_0489_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][0] ),
    .CLK(_0146_));
 sg13g2_dfrbpq_1 _5062_ (.RESET_B(net59),
    .D(_0490_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][1] ),
    .CLK(_0147_));
 sg13g2_dfrbpq_1 _5063_ (.RESET_B(net55),
    .D(_0491_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][2] ),
    .CLK(_0148_));
 sg13g2_dfrbpq_1 _5064_ (.RESET_B(net262),
    .D(_0492_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[3][3] ),
    .CLK(_0149_));
 sg13g2_dfrbpq_1 _5065_ (.RESET_B(net263),
    .D(_0002_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[0] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _5066_ (.RESET_B(net264),
    .D(_0003_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[1] ),
    .CLK(net635));
 sg13g2_dfrbpq_2 _5067_ (.RESET_B(net402),
    .D(_0000_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[2] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _5068_ (.RESET_B(net51),
    .D(_0001_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.state[3] ),
    .CLK(net635));
 sg13g2_dfrbpq_1 _5069_ (.RESET_B(net47),
    .D(_0493_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][0] ),
    .CLK(_0150_));
 sg13g2_dfrbpq_1 _5070_ (.RESET_B(net43),
    .D(_0494_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][1] ),
    .CLK(_0151_));
 sg13g2_dfrbpq_1 _5071_ (.RESET_B(net39),
    .D(_0495_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][2] ),
    .CLK(_0152_));
 sg13g2_dfrbpq_1 _5072_ (.RESET_B(net35),
    .D(_0496_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[15][3] ),
    .CLK(_0153_));
 sg13g2_dfrbpq_1 _5073_ (.RESET_B(net31),
    .D(_0497_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][0] ),
    .CLK(_0154_));
 sg13g2_dfrbpq_1 _5074_ (.RESET_B(net399),
    .D(_0498_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][1] ),
    .CLK(_0155_));
 sg13g2_dfrbpq_1 _5075_ (.RESET_B(net395),
    .D(_0499_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][2] ),
    .CLK(_0156_));
 sg13g2_dfrbpq_1 _5076_ (.RESET_B(net391),
    .D(_0500_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[11][3] ),
    .CLK(_0157_));
 sg13g2_dfrbpq_1 _5077_ (.RESET_B(net387),
    .D(_0501_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][0] ),
    .CLK(_0158_));
 sg13g2_dfrbpq_1 _5078_ (.RESET_B(net383),
    .D(_0502_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][1] ),
    .CLK(_0159_));
 sg13g2_dfrbpq_1 _5079_ (.RESET_B(net379),
    .D(_0503_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][2] ),
    .CLK(_0160_));
 sg13g2_dfrbpq_1 _5080_ (.RESET_B(net375),
    .D(_0504_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[13][3] ),
    .CLK(_0161_));
 sg13g2_dfrbpq_1 _5081_ (.RESET_B(net371),
    .D(_0505_),
    .Q(\green_tmds_par[2] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _5082_ (.RESET_B(net369),
    .D(_0506_),
    .Q(\green_tmds_par[6] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _5083_ (.RESET_B(net367),
    .D(_0507_),
    .Q(\green_tmds_par[8] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5084_ (.RESET_B(net365),
    .D(_0508_),
    .Q(\green_tmds_par[9] ),
    .CLK(net646));
 sg13g2_dfrbpq_1 _5085_ (.RESET_B(net363),
    .D(_0509_),
    .Q(\tmds_red.dc_balancing_reg[0] ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _5086_ (.RESET_B(net361),
    .D(_0510_),
    .Q(\tmds_red.dc_balancing_reg[1] ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _5087_ (.RESET_B(net359),
    .D(_0511_),
    .Q(\tmds_red.dc_balancing_reg[2] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _5088_ (.RESET_B(net357),
    .D(_0512_),
    .Q(\tmds_red.dc_balancing_reg[3] ),
    .CLK(net644));
 sg13g2_dfrbpq_2 _5089_ (.RESET_B(net355),
    .D(_0513_),
    .Q(\tmds_red.dc_balancing_reg[4] ),
    .CLK(net644));
 sg13g2_dfrbpq_1 _5090_ (.RESET_B(net353),
    .D(_0514_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][0] ),
    .CLK(_0162_));
 sg13g2_dfrbpq_1 _5091_ (.RESET_B(net349),
    .D(_0515_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][1] ),
    .CLK(_0163_));
 sg13g2_dfrbpq_1 _5092_ (.RESET_B(net322),
    .D(_0516_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][2] ),
    .CLK(_0164_));
 sg13g2_dfrbpq_1 _5093_ (.RESET_B(net318),
    .D(_0517_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[37][3] ),
    .CLK(_0165_));
 sg13g2_dfrbpq_1 _5094_ (.RESET_B(net314),
    .D(_0518_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][0] ),
    .CLK(_0166_));
 sg13g2_dfrbpq_1 _5095_ (.RESET_B(net310),
    .D(_0519_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][1] ),
    .CLK(_0167_));
 sg13g2_dfrbpq_1 _5096_ (.RESET_B(net306),
    .D(_0520_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][2] ),
    .CLK(_0168_));
 sg13g2_dfrbpq_1 _5097_ (.RESET_B(net302),
    .D(_0521_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[36][3] ),
    .CLK(_0169_));
 sg13g2_dfrbpq_1 _5098_ (.RESET_B(net299),
    .D(_0522_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][0] ),
    .CLK(_0170_));
 sg13g2_dfrbpq_1 _5099_ (.RESET_B(net295),
    .D(_0523_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][1] ),
    .CLK(_0171_));
 sg13g2_dfrbpq_1 _5100_ (.RESET_B(net291),
    .D(_0524_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][2] ),
    .CLK(_0172_));
 sg13g2_dfrbpq_1 _5101_ (.RESET_B(net287),
    .D(_0525_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[35][3] ),
    .CLK(_0173_));
 sg13g2_dfrbpq_1 _5102_ (.RESET_B(net283),
    .D(_0526_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][0] ),
    .CLK(_0174_));
 sg13g2_dfrbpq_1 _5103_ (.RESET_B(net279),
    .D(_0527_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][1] ),
    .CLK(_0175_));
 sg13g2_dfrbpq_1 _5104_ (.RESET_B(net275),
    .D(_0528_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][2] ),
    .CLK(_0176_));
 sg13g2_dfrbpq_1 _5105_ (.RESET_B(net271),
    .D(_0529_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[34][3] ),
    .CLK(_0177_));
 sg13g2_dfrbpq_1 _5106_ (.RESET_B(net268),
    .D(_0530_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][0] ),
    .CLK(_0178_));
 sg13g2_dfrbpq_1 _5107_ (.RESET_B(net260),
    .D(_0531_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][1] ),
    .CLK(_0179_));
 sg13g2_dfrbpq_1 _5108_ (.RESET_B(net256),
    .D(_0532_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][2] ),
    .CLK(_0180_));
 sg13g2_dfrbpq_1 _5109_ (.RESET_B(net252),
    .D(_0533_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[33][3] ),
    .CLK(_0181_));
 sg13g2_dfrbpq_1 _5110_ (.RESET_B(net248),
    .D(_0534_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][0] ),
    .CLK(_0182_));
 sg13g2_dfrbpq_1 _5111_ (.RESET_B(net244),
    .D(_0535_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][1] ),
    .CLK(_0183_));
 sg13g2_dfrbpq_1 _5112_ (.RESET_B(net240),
    .D(_0536_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][2] ),
    .CLK(_0184_));
 sg13g2_dfrbpq_1 _5113_ (.RESET_B(net236),
    .D(_0537_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[32][3] ),
    .CLK(_0185_));
 sg13g2_dfrbpq_1 _5114_ (.RESET_B(net233),
    .D(_0538_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][0] ),
    .CLK(_0186_));
 sg13g2_dfrbpq_1 _5115_ (.RESET_B(net229),
    .D(_0539_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][1] ),
    .CLK(_0187_));
 sg13g2_dfrbpq_1 _5116_ (.RESET_B(net225),
    .D(_0540_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][2] ),
    .CLK(_0188_));
 sg13g2_dfrbpq_1 _5117_ (.RESET_B(net221),
    .D(_0541_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[31][3] ),
    .CLK(_0189_));
 sg13g2_dfrbpq_1 _5118_ (.RESET_B(net217),
    .D(_0542_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][0] ),
    .CLK(_0190_));
 sg13g2_dfrbpq_1 _5119_ (.RESET_B(net213),
    .D(_0543_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][1] ),
    .CLK(_0191_));
 sg13g2_dfrbpq_1 _5120_ (.RESET_B(net209),
    .D(_0544_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][2] ),
    .CLK(_0192_));
 sg13g2_dfrbpq_1 _5121_ (.RESET_B(net205),
    .D(_0545_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[30][3] ),
    .CLK(_0193_));
 sg13g2_dfrbpq_1 _5122_ (.RESET_B(net201),
    .D(_0546_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][0] ),
    .CLK(_0194_));
 sg13g2_dfrbpq_1 _5123_ (.RESET_B(net197),
    .D(_0547_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][1] ),
    .CLK(_0195_));
 sg13g2_dfrbpq_1 _5124_ (.RESET_B(net193),
    .D(_0548_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][2] ),
    .CLK(_0196_));
 sg13g2_dfrbpq_1 _5125_ (.RESET_B(net189),
    .D(_0549_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[2][3] ),
    .CLK(_0197_));
 sg13g2_dfrbpq_1 _5126_ (.RESET_B(net185),
    .D(_0550_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][0] ),
    .CLK(_0198_));
 sg13g2_dfrbpq_1 _5127_ (.RESET_B(net181),
    .D(_0551_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][1] ),
    .CLK(_0199_));
 sg13g2_dfrbpq_1 _5128_ (.RESET_B(net177),
    .D(_0552_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][2] ),
    .CLK(_0200_));
 sg13g2_dfrbpq_1 _5129_ (.RESET_B(net173),
    .D(_0553_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[28][3] ),
    .CLK(_0201_));
 sg13g2_dfrbpq_1 _5130_ (.RESET_B(net169),
    .D(_0554_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][0] ),
    .CLK(_0202_));
 sg13g2_dfrbpq_1 _5131_ (.RESET_B(net165),
    .D(_0555_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][1] ),
    .CLK(_0203_));
 sg13g2_dfrbpq_1 _5132_ (.RESET_B(net161),
    .D(_0556_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][2] ),
    .CLK(_0204_));
 sg13g2_dfrbpq_1 _5133_ (.RESET_B(net152),
    .D(_0557_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[27][3] ),
    .CLK(_0205_));
 sg13g2_dfrbpq_1 _5134_ (.RESET_B(net136),
    .D(_0558_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][0] ),
    .CLK(_0206_));
 sg13g2_dfrbpq_1 _5135_ (.RESET_B(net128),
    .D(_0559_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][1] ),
    .CLK(_0207_));
 sg13g2_dfrbpq_1 _5136_ (.RESET_B(net120),
    .D(_0560_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][2] ),
    .CLK(_0208_));
 sg13g2_dfrbpq_1 _5137_ (.RESET_B(net112),
    .D(_0561_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[26][3] ),
    .CLK(_0209_));
 sg13g2_dfrbpq_1 _5138_ (.RESET_B(net104),
    .D(_0562_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][0] ),
    .CLK(_0210_));
 sg13g2_dfrbpq_1 _5139_ (.RESET_B(net86),
    .D(_0563_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][1] ),
    .CLK(_0211_));
 sg13g2_dfrbpq_1 _5140_ (.RESET_B(net78),
    .D(_0564_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][2] ),
    .CLK(_0212_));
 sg13g2_dfrbpq_1 _5141_ (.RESET_B(net69),
    .D(_0565_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[25][3] ),
    .CLK(_0213_));
 sg13g2_dfrbpq_1 _5142_ (.RESET_B(net61),
    .D(_0566_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][0] ),
    .CLK(_0214_));
 sg13g2_dfrbpq_1 _5143_ (.RESET_B(net53),
    .D(_0567_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][1] ),
    .CLK(_0215_));
 sg13g2_dfrbpq_1 _5144_ (.RESET_B(net45),
    .D(_0568_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][2] ),
    .CLK(_0216_));
 sg13g2_dfrbpq_1 _5145_ (.RESET_B(net37),
    .D(_0569_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[24][3] ),
    .CLK(_0217_));
 sg13g2_dfrbpq_1 _5146_ (.RESET_B(net401),
    .D(_0570_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][0] ),
    .CLK(_0218_));
 sg13g2_dfrbpq_1 _5147_ (.RESET_B(net393),
    .D(_0571_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][1] ),
    .CLK(_0219_));
 sg13g2_dfrbpq_1 _5148_ (.RESET_B(net385),
    .D(_0572_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][2] ),
    .CLK(_0220_));
 sg13g2_dfrbpq_1 _5149_ (.RESET_B(net377),
    .D(_0573_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[23][3] ),
    .CLK(_0221_));
 sg13g2_dfrbpq_1 _5150_ (.RESET_B(net351),
    .D(_0574_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][0] ),
    .CLK(_0222_));
 sg13g2_dfrbpq_1 _5151_ (.RESET_B(net320),
    .D(_0575_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][1] ),
    .CLK(_0223_));
 sg13g2_dfrbpq_1 _5152_ (.RESET_B(net312),
    .D(_0576_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][2] ),
    .CLK(_0224_));
 sg13g2_dfrbpq_1 _5153_ (.RESET_B(net304),
    .D(_0577_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[22][3] ),
    .CLK(_0225_));
 sg13g2_dfrbpq_1 _5154_ (.RESET_B(net297),
    .D(_0578_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][0] ),
    .CLK(_0226_));
 sg13g2_dfrbpq_1 _5155_ (.RESET_B(net289),
    .D(_0579_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][1] ),
    .CLK(_0227_));
 sg13g2_dfrbpq_1 _5156_ (.RESET_B(net281),
    .D(_0580_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][2] ),
    .CLK(_0228_));
 sg13g2_dfrbpq_1 _5157_ (.RESET_B(net273),
    .D(_0581_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[21][3] ),
    .CLK(_0229_));
 sg13g2_dfrbpq_1 _5158_ (.RESET_B(net266),
    .D(_0582_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][0] ),
    .CLK(_0230_));
 sg13g2_dfrbpq_1 _5159_ (.RESET_B(net254),
    .D(_0583_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][1] ),
    .CLK(_0231_));
 sg13g2_dfrbpq_1 _5160_ (.RESET_B(net246),
    .D(_0584_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][2] ),
    .CLK(_0232_));
 sg13g2_dfrbpq_1 _5161_ (.RESET_B(net238),
    .D(_0585_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[20][3] ),
    .CLK(_0233_));
 sg13g2_dfrbpq_1 _5162_ (.RESET_B(net231),
    .D(_0586_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][0] ),
    .CLK(_0234_));
 sg13g2_dfrbpq_1 _5163_ (.RESET_B(net223),
    .D(_0587_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][1] ),
    .CLK(_0235_));
 sg13g2_dfrbpq_1 _5164_ (.RESET_B(net215),
    .D(_0588_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][2] ),
    .CLK(_0236_));
 sg13g2_dfrbpq_1 _5165_ (.RESET_B(net207),
    .D(_0589_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[1][3] ),
    .CLK(_0237_));
 sg13g2_dfrbpq_1 _5166_ (.RESET_B(net199),
    .D(_0590_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][0] ),
    .CLK(_0238_));
 sg13g2_dfrbpq_1 _5167_ (.RESET_B(net191),
    .D(_0591_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][1] ),
    .CLK(_0239_));
 sg13g2_dfrbpq_1 _5168_ (.RESET_B(net183),
    .D(_0592_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][2] ),
    .CLK(_0240_));
 sg13g2_dfrbpq_1 _5169_ (.RESET_B(net175),
    .D(_0593_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[18][3] ),
    .CLK(_0241_));
 sg13g2_dfrbpq_1 _5170_ (.RESET_B(net167),
    .D(_0594_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][0] ),
    .CLK(_0242_));
 sg13g2_dfrbpq_1 _5171_ (.RESET_B(net159),
    .D(_0595_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][1] ),
    .CLK(_0243_));
 sg13g2_dfrbpq_1 _5172_ (.RESET_B(net132),
    .D(_0596_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][2] ),
    .CLK(_0244_));
 sg13g2_dfrbpq_1 _5173_ (.RESET_B(net116),
    .D(_0597_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[17][3] ),
    .CLK(_0245_));
 sg13g2_dfrbpq_1 _5174_ (.RESET_B(net100),
    .D(_0598_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][0] ),
    .CLK(_0246_));
 sg13g2_dfrbpq_1 _5175_ (.RESET_B(net74),
    .D(_0599_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][1] ),
    .CLK(_0247_));
 sg13g2_dfrbpq_1 _5176_ (.RESET_B(net57),
    .D(_0600_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][2] ),
    .CLK(_0248_));
 sg13g2_dfrbpq_1 _5177_ (.RESET_B(net41),
    .D(_0601_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[16][3] ),
    .CLK(_0249_));
 sg13g2_dfrbpq_1 _5178_ (.RESET_B(net397),
    .D(_0602_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][0] ),
    .CLK(_0250_));
 sg13g2_dfrbpq_1 _5179_ (.RESET_B(net381),
    .D(_0603_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][1] ),
    .CLK(_0251_));
 sg13g2_dfrbpq_1 _5180_ (.RESET_B(net347),
    .D(_0604_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][2] ),
    .CLK(_0252_));
 sg13g2_dfrbpq_1 _5181_ (.RESET_B(net308),
    .D(_0605_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[7][3] ),
    .CLK(_0253_));
 sg13g2_dfrbpq_1 _5182_ (.RESET_B(net293),
    .D(_0606_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][0] ),
    .CLK(_0254_));
 sg13g2_dfrbpq_1 _5183_ (.RESET_B(net277),
    .D(_0607_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][1] ),
    .CLK(_0255_));
 sg13g2_dfrbpq_1 _5184_ (.RESET_B(net258),
    .D(_0608_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][2] ),
    .CLK(_0256_));
 sg13g2_dfrbpq_1 _5185_ (.RESET_B(net242),
    .D(_0609_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[10][3] ),
    .CLK(_0257_));
 sg13g2_dfrbpq_1 _5186_ (.RESET_B(net227),
    .D(_0610_),
    .Q(\blue_tmds_par[0] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5187_ (.RESET_B(net219),
    .D(_0611_),
    .Q(\blue_tmds_par[1] ),
    .CLK(net643));
 sg13g2_dfrbpq_1 _5188_ (.RESET_B(net211),
    .D(_0612_),
    .Q(\blue_tmds_par[2] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5189_ (.RESET_B(net203),
    .D(_0613_),
    .Q(\blue_tmds_par[3] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5190_ (.RESET_B(net195),
    .D(_0614_),
    .Q(\blue_tmds_par[5] ),
    .CLK(net638));
 sg13g2_dfrbpq_1 _5191_ (.RESET_B(net187),
    .D(_0615_),
    .Q(\blue_tmds_par[6] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5192_ (.RESET_B(net179),
    .D(_0616_),
    .Q(\blue_tmds_par[7] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5193_ (.RESET_B(net171),
    .D(_0617_),
    .Q(\blue_tmds_par[8] ),
    .CLK(net637));
 sg13g2_dfrbpq_1 _5194_ (.RESET_B(net163),
    .D(_0618_),
    .Q(\blue_tmds_par[9] ),
    .CLK(net637));
 sg13g2_dfrbpq_2 _5195_ (.RESET_B(net148),
    .D(_0619_),
    .Q(\tmds_green.dc_balancing_reg[1] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _5196_ (.RESET_B(net124),
    .D(_0620_),
    .Q(\tmds_green.dc_balancing_reg[2] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _5197_ (.RESET_B(net108),
    .D(_0621_),
    .Q(\tmds_green.dc_balancing_reg[3] ),
    .CLK(net645));
 sg13g2_dfrbpq_2 _5198_ (.RESET_B(net82),
    .D(_0622_),
    .Q(\tmds_green.dc_balancing_reg[4] ),
    .CLK(net645));
 sg13g2_dfrbpq_1 _5199_ (.RESET_B(net65),
    .D(net407),
    .Q(\clockdiv.q0 ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _5200_ (.RESET_B(net49),
    .D(_0624_),
    .Q(\tmds_blue.dc_balancing_reg[1] ),
    .CLK(net639));
 sg13g2_dfrbpq_1 _5201_ (.RESET_B(net33),
    .D(_0625_),
    .Q(\tmds_blue.dc_balancing_reg[2] ),
    .CLK(net639));
 sg13g2_dfrbpq_2 _5202_ (.RESET_B(net389),
    .D(_0626_),
    .Q(\tmds_blue.dc_balancing_reg[3] ),
    .CLK(net638));
 sg13g2_dfrbpq_2 _5203_ (.RESET_B(net373),
    .D(_0627_),
    .Q(\tmds_blue.dc_balancing_reg[4] ),
    .CLK(net638));
 sg13g2_dfrbpq_1 _5204_ (.RESET_B(net316),
    .D(_0628_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][0] ),
    .CLK(_0258_));
 sg13g2_dfrbpq_1 _5205_ (.RESET_B(net285),
    .D(_0629_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][1] ),
    .CLK(_0259_));
 sg13g2_dfrbpq_1 _5206_ (.RESET_B(net250),
    .D(_0630_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][2] ),
    .CLK(_0260_));
 sg13g2_dfrbpq_1 _5207_ (.RESET_B(net403),
    .D(_0631_),
    .Q(\videogen.test_lut_thingy.pixel_feeder_inst.row[14][3] ),
    .CLK(_0261_));
 sg13g2_dfrbpq_1 _5208_ (.RESET_B(net803),
    .D(\serialize.n428[0] ),
    .Q(\serialize.n453 ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5209_ (.RESET_B(net803),
    .D(\serialize.n428[1] ),
    .Q(\serialize.n455 ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5210_ (.RESET_B(net802),
    .D(\serialize.n428[2] ),
    .Q(\serialize.n414[0] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5211_ (.RESET_B(net803),
    .D(\serialize.n428[3] ),
    .Q(\serialize.n414[1] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5212_ (.RESET_B(net802),
    .D(\serialize.n428[4] ),
    .Q(\serialize.n414[2] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5213_ (.RESET_B(net803),
    .D(\serialize.n428[5] ),
    .Q(\serialize.n414[3] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5214_ (.RESET_B(net801),
    .D(\serialize.n428[6] ),
    .Q(\serialize.n414[4] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5215_ (.RESET_B(net803),
    .D(\serialize.n428[7] ),
    .Q(\serialize.n414[5] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5216_ (.RESET_B(net801),
    .D(\serialize.n428[8] ),
    .Q(\serialize.n414[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5217_ (.RESET_B(net804),
    .D(\serialize.n428[9] ),
    .Q(\serialize.n414[7] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5218_ (.RESET_B(net803),
    .D(\serialize.n431[0] ),
    .Q(\serialize.n459 ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5219_ (.RESET_B(net803),
    .D(\serialize.n431[1] ),
    .Q(\serialize.n461 ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5220_ (.RESET_B(net805),
    .D(\serialize.n431[2] ),
    .Q(\serialize.n420[0] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5221_ (.RESET_B(net804),
    .D(\serialize.n431[3] ),
    .Q(\serialize.n420[1] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5222_ (.RESET_B(net804),
    .D(\serialize.n431[4] ),
    .Q(\serialize.n420[2] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5223_ (.RESET_B(net804),
    .D(\serialize.n431[5] ),
    .Q(\serialize.n420[3] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5224_ (.RESET_B(net804),
    .D(net420),
    .Q(\serialize.n420[4] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5225_ (.RESET_B(net800),
    .D(net694),
    .Q(\serialize.n420[6] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5226_ (.RESET_B(net804),
    .D(\serialize.n429[0] ),
    .Q(\serialize.n456 ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5227_ (.RESET_B(net804),
    .D(\serialize.n429[1] ),
    .Q(\serialize.n458 ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5228_ (.RESET_B(net799),
    .D(\serialize.n429[2] ),
    .Q(\serialize.n417[0] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5229_ (.RESET_B(net799),
    .D(net434),
    .Q(\serialize.n417[1] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5230_ (.RESET_B(net800),
    .D(net444),
    .Q(\serialize.n417[2] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5231_ (.RESET_B(net800),
    .D(\serialize.n429[5] ),
    .Q(\serialize.n417[3] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5232_ (.RESET_B(net800),
    .D(\serialize.n429[6] ),
    .Q(\serialize.n417[4] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5233_ (.RESET_B(net799),
    .D(\serialize.n429[7] ),
    .Q(\serialize.n417[5] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5234_ (.RESET_B(net799),
    .D(\serialize.n429[8] ),
    .Q(\serialize.n417[6] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5235_ (.RESET_B(net799),
    .D(\serialize.n429[9] ),
    .Q(\serialize.n417[7] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _5236_ (.RESET_B(net801),
    .D(\serialize.n433[0] ),
    .Q(\serialize.bit_cnt[0] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5237_ (.RESET_B(net801),
    .D(\serialize.n433[1] ),
    .Q(\serialize.bit_cnt[1] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5238_ (.RESET_B(net801),
    .D(net416),
    .Q(_0004_),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5239_ (.RESET_B(net805),
    .D(\serialize.n427[0] ),
    .Q(\serialize.n450 ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5240_ (.RESET_B(net805),
    .D(\serialize.n427[1] ),
    .Q(\serialize.n452 ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5241_ (.RESET_B(net802),
    .D(\serialize.n427[2] ),
    .Q(\serialize.n411[0] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5242_ (.RESET_B(net802),
    .D(\serialize.n427[3] ),
    .Q(\serialize.n411[1] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5243_ (.RESET_B(net802),
    .D(\serialize.n427[4] ),
    .Q(\serialize.n411[2] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5244_ (.RESET_B(net805),
    .D(\serialize.n427[5] ),
    .Q(\serialize.n411[3] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5245_ (.RESET_B(net802),
    .D(\serialize.n427[6] ),
    .Q(\serialize.n411[4] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5246_ (.RESET_B(net802),
    .D(\serialize.n427[7] ),
    .Q(\serialize.n411[5] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5247_ (.RESET_B(net801),
    .D(\serialize.n427[8] ),
    .Q(\serialize.n411[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _5248_ (.RESET_B(net802),
    .D(\serialize.n427[9] ),
    .Q(\serialize.n411[7] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_tiehi _4909__32 (.L_HI(net32));
 sg13g2_tiehi _5201__33 (.L_HI(net33));
 sg13g2_tiehi _4908__34 (.L_HI(net34));
 sg13g2_tiehi _5072__35 (.L_HI(net35));
 sg13g2_tiehi _4907__36 (.L_HI(net36));
 sg13g2_tiehi _5145__37 (.L_HI(net37));
 sg13g2_tiehi _4906__38 (.L_HI(net38));
 sg13g2_tiehi _5071__39 (.L_HI(net39));
 sg13g2_tiehi _4905__40 (.L_HI(net40));
 sg13g2_tiehi _5177__41 (.L_HI(net41));
 sg13g2_tiehi _4904__42 (.L_HI(net42));
 sg13g2_tiehi _5070__43 (.L_HI(net43));
 sg13g2_tiehi _4903__44 (.L_HI(net44));
 sg13g2_tiehi _5144__45 (.L_HI(net45));
 sg13g2_tiehi _4902__46 (.L_HI(net46));
 sg13g2_tiehi _5069__47 (.L_HI(net47));
 sg13g2_tiehi _4901__48 (.L_HI(net48));
 sg13g2_tiehi _5200__49 (.L_HI(net49));
 sg13g2_tiehi _4900__50 (.L_HI(net50));
 sg13g2_tiehi _5068__51 (.L_HI(net51));
 sg13g2_tiehi _4899__52 (.L_HI(net52));
 sg13g2_tiehi _5143__53 (.L_HI(net53));
 sg13g2_tiehi _4898__54 (.L_HI(net54));
 sg13g2_tiehi _5063__55 (.L_HI(net55));
 sg13g2_tiehi _4897__56 (.L_HI(net56));
 sg13g2_tiehi _5176__57 (.L_HI(net57));
 sg13g2_tiehi _4896__58 (.L_HI(net58));
 sg13g2_tiehi _5062__59 (.L_HI(net59));
 sg13g2_tiehi _4895__60 (.L_HI(net60));
 sg13g2_tiehi _5142__61 (.L_HI(net61));
 sg13g2_tiehi _4894__62 (.L_HI(net62));
 sg13g2_tiehi _5061__63 (.L_HI(net63));
 sg13g2_tiehi _4893__64 (.L_HI(net64));
 sg13g2_tiehi _5199__65 (.L_HI(net65));
 sg13g2_tiehi _4892__66 (.L_HI(net66));
 sg13g2_tiehi _5060__67 (.L_HI(net67));
 sg13g2_tiehi _4891__68 (.L_HI(net68));
 sg13g2_tiehi _5141__69 (.L_HI(net69));
 sg13g2_tiehi _4890__70 (.L_HI(net70));
 sg13g2_tiehi _4889__71 (.L_HI(net71));
 sg13g2_tiehi _5059__72 (.L_HI(net72));
 sg13g2_tiehi _4888__73 (.L_HI(net73));
 sg13g2_tiehi _5175__74 (.L_HI(net74));
 sg13g2_tiehi _4887__75 (.L_HI(net75));
 sg13g2_tiehi _5058__76 (.L_HI(net76));
 sg13g2_tiehi _4886__77 (.L_HI(net77));
 sg13g2_tiehi _5140__78 (.L_HI(net78));
 sg13g2_tiehi _4885__79 (.L_HI(net79));
 sg13g2_tiehi _5057__80 (.L_HI(net80));
 sg13g2_tiehi _4884__81 (.L_HI(net81));
 sg13g2_tiehi _5198__82 (.L_HI(net82));
 sg13g2_tiehi _4883__83 (.L_HI(net83));
 sg13g2_tiehi _5056__84 (.L_HI(net84));
 sg13g2_tiehi _4882__85 (.L_HI(net85));
 sg13g2_tiehi _5139__86 (.L_HI(net86));
 sg13g2_tiehi _4881__87 (.L_HI(net87));
 sg13g2_tiehi _4880__88 (.L_HI(net88));
 sg13g2_tiehi _4879__89 (.L_HI(net89));
 sg13g2_tiehi _4878__90 (.L_HI(net90));
 sg13g2_tiehi _4877__91 (.L_HI(net91));
 sg13g2_tiehi _4876__92 (.L_HI(net92));
 sg13g2_tiehi _4875__93 (.L_HI(net93));
 sg13g2_tiehi _4874__94 (.L_HI(net94));
 sg13g2_tiehi _4873__95 (.L_HI(net95));
 sg13g2_tiehi _4872__96 (.L_HI(net96));
 sg13g2_tiehi _4871__97 (.L_HI(net97));
 sg13g2_tiehi _5055__98 (.L_HI(net98));
 sg13g2_tiehi _4870__99 (.L_HI(net99));
 sg13g2_tiehi _5174__100 (.L_HI(net100));
 sg13g2_tiehi _4869__101 (.L_HI(net101));
 sg13g2_tiehi _5054__102 (.L_HI(net102));
 sg13g2_tiehi _4868__103 (.L_HI(net103));
 sg13g2_tiehi _5138__104 (.L_HI(net104));
 sg13g2_tiehi _4867__105 (.L_HI(net105));
 sg13g2_tiehi _5053__106 (.L_HI(net106));
 sg13g2_tiehi _4866__107 (.L_HI(net107));
 sg13g2_tiehi _5197__108 (.L_HI(net108));
 sg13g2_tiehi _4865__109 (.L_HI(net109));
 sg13g2_tiehi _5052__110 (.L_HI(net110));
 sg13g2_tiehi _4864__111 (.L_HI(net111));
 sg13g2_tiehi _5137__112 (.L_HI(net112));
 sg13g2_tiehi _4863__113 (.L_HI(net113));
 sg13g2_tiehi _5051__114 (.L_HI(net114));
 sg13g2_tiehi _4862__115 (.L_HI(net115));
 sg13g2_tiehi _5173__116 (.L_HI(net116));
 sg13g2_tiehi _4861__117 (.L_HI(net117));
 sg13g2_tiehi _5050__118 (.L_HI(net118));
 sg13g2_tiehi _4860__119 (.L_HI(net119));
 sg13g2_tiehi _5136__120 (.L_HI(net120));
 sg13g2_tiehi _4859__121 (.L_HI(net121));
 sg13g2_tiehi _5049__122 (.L_HI(net122));
 sg13g2_tiehi _4858__123 (.L_HI(net123));
 sg13g2_tiehi _5196__124 (.L_HI(net124));
 sg13g2_tiehi _4857__125 (.L_HI(net125));
 sg13g2_tiehi _5048__126 (.L_HI(net126));
 sg13g2_tiehi _4856__127 (.L_HI(net127));
 sg13g2_tiehi _5135__128 (.L_HI(net128));
 sg13g2_tiehi _4855__129 (.L_HI(net129));
 sg13g2_tiehi _5047__130 (.L_HI(net130));
 sg13g2_tiehi _4854__131 (.L_HI(net131));
 sg13g2_tiehi _5172__132 (.L_HI(net132));
 sg13g2_tiehi _4853__133 (.L_HI(net133));
 sg13g2_tiehi _5046__134 (.L_HI(net134));
 sg13g2_tiehi _4852__135 (.L_HI(net135));
 sg13g2_tiehi _5134__136 (.L_HI(net136));
 sg13g2_tiehi _4851__137 (.L_HI(net137));
 sg13g2_tiehi _4850__138 (.L_HI(net138));
 sg13g2_tiehi _4849__139 (.L_HI(net139));
 sg13g2_tiehi _4848__140 (.L_HI(net140));
 sg13g2_tiehi _4847__141 (.L_HI(net141));
 sg13g2_tiehi _4846__142 (.L_HI(net142));
 sg13g2_tiehi _4845__143 (.L_HI(net143));
 sg13g2_tiehi _4844__144 (.L_HI(net144));
 sg13g2_tiehi _4843__145 (.L_HI(net145));
 sg13g2_tiehi _5045__146 (.L_HI(net146));
 sg13g2_tiehi _4842__147 (.L_HI(net147));
 sg13g2_tiehi _5195__148 (.L_HI(net148));
 sg13g2_tiehi _4841__149 (.L_HI(net149));
 sg13g2_tiehi _5044__150 (.L_HI(net150));
 sg13g2_tiehi _4840__151 (.L_HI(net151));
 sg13g2_tiehi _5133__152 (.L_HI(net152));
 sg13g2_tiehi _4839__153 (.L_HI(net153));
 sg13g2_tiehi _4838__154 (.L_HI(net154));
 sg13g2_tiehi _4837__155 (.L_HI(net155));
 sg13g2_tiehi _4836__156 (.L_HI(net156));
 sg13g2_tiehi _5043__157 (.L_HI(net157));
 sg13g2_tiehi _4835__158 (.L_HI(net158));
 sg13g2_tiehi _5171__159 (.L_HI(net159));
 sg13g2_tiehi _5042__160 (.L_HI(net160));
 sg13g2_tiehi _5132__161 (.L_HI(net161));
 sg13g2_tiehi _5041__162 (.L_HI(net162));
 sg13g2_tiehi _5194__163 (.L_HI(net163));
 sg13g2_tiehi _5040__164 (.L_HI(net164));
 sg13g2_tiehi _5131__165 (.L_HI(net165));
 sg13g2_tiehi _5039__166 (.L_HI(net166));
 sg13g2_tiehi _5170__167 (.L_HI(net167));
 sg13g2_tiehi _5038__168 (.L_HI(net168));
 sg13g2_tiehi _5130__169 (.L_HI(net169));
 sg13g2_tiehi _5037__170 (.L_HI(net170));
 sg13g2_tiehi _5193__171 (.L_HI(net171));
 sg13g2_tiehi _5036__172 (.L_HI(net172));
 sg13g2_tiehi _5129__173 (.L_HI(net173));
 sg13g2_tiehi _5035__174 (.L_HI(net174));
 sg13g2_tiehi _5169__175 (.L_HI(net175));
 sg13g2_tiehi _5034__176 (.L_HI(net176));
 sg13g2_tiehi _5128__177 (.L_HI(net177));
 sg13g2_tiehi _5033__178 (.L_HI(net178));
 sg13g2_tiehi _5192__179 (.L_HI(net179));
 sg13g2_tiehi _5032__180 (.L_HI(net180));
 sg13g2_tiehi _5127__181 (.L_HI(net181));
 sg13g2_tiehi _5031__182 (.L_HI(net182));
 sg13g2_tiehi _5168__183 (.L_HI(net183));
 sg13g2_tiehi _5030__184 (.L_HI(net184));
 sg13g2_tiehi _5126__185 (.L_HI(net185));
 sg13g2_tiehi _5029__186 (.L_HI(net186));
 sg13g2_tiehi _5191__187 (.L_HI(net187));
 sg13g2_tiehi _5028__188 (.L_HI(net188));
 sg13g2_tiehi _5125__189 (.L_HI(net189));
 sg13g2_tiehi _5027__190 (.L_HI(net190));
 sg13g2_tiehi _5167__191 (.L_HI(net191));
 sg13g2_tiehi _5026__192 (.L_HI(net192));
 sg13g2_tiehi _5124__193 (.L_HI(net193));
 sg13g2_tiehi _5025__194 (.L_HI(net194));
 sg13g2_tiehi _5190__195 (.L_HI(net195));
 sg13g2_tiehi _5024__196 (.L_HI(net196));
 sg13g2_tiehi _5123__197 (.L_HI(net197));
 sg13g2_tiehi _5023__198 (.L_HI(net198));
 sg13g2_tiehi _5166__199 (.L_HI(net199));
 sg13g2_tiehi _5022__200 (.L_HI(net200));
 sg13g2_tiehi _5122__201 (.L_HI(net201));
 sg13g2_tiehi _5021__202 (.L_HI(net202));
 sg13g2_tiehi _5189__203 (.L_HI(net203));
 sg13g2_tiehi _5020__204 (.L_HI(net204));
 sg13g2_tiehi _5121__205 (.L_HI(net205));
 sg13g2_tiehi _5019__206 (.L_HI(net206));
 sg13g2_tiehi _5165__207 (.L_HI(net207));
 sg13g2_tiehi _5018__208 (.L_HI(net208));
 sg13g2_tiehi _5120__209 (.L_HI(net209));
 sg13g2_tiehi _5017__210 (.L_HI(net210));
 sg13g2_tiehi _5188__211 (.L_HI(net211));
 sg13g2_tiehi _5016__212 (.L_HI(net212));
 sg13g2_tiehi _5119__213 (.L_HI(net213));
 sg13g2_tiehi _5015__214 (.L_HI(net214));
 sg13g2_tiehi _5164__215 (.L_HI(net215));
 sg13g2_tiehi _5014__216 (.L_HI(net216));
 sg13g2_tiehi _5118__217 (.L_HI(net217));
 sg13g2_tiehi _5013__218 (.L_HI(net218));
 sg13g2_tiehi _5187__219 (.L_HI(net219));
 sg13g2_tiehi _5012__220 (.L_HI(net220));
 sg13g2_tiehi _5117__221 (.L_HI(net221));
 sg13g2_tiehi _5011__222 (.L_HI(net222));
 sg13g2_tiehi _5163__223 (.L_HI(net223));
 sg13g2_tiehi _5010__224 (.L_HI(net224));
 sg13g2_tiehi _5116__225 (.L_HI(net225));
 sg13g2_tiehi _5009__226 (.L_HI(net226));
 sg13g2_tiehi _5186__227 (.L_HI(net227));
 sg13g2_tiehi _5008__228 (.L_HI(net228));
 sg13g2_tiehi _5115__229 (.L_HI(net229));
 sg13g2_tiehi _5007__230 (.L_HI(net230));
 sg13g2_tiehi _5162__231 (.L_HI(net231));
 sg13g2_tiehi _5006__232 (.L_HI(net232));
 sg13g2_tiehi _5114__233 (.L_HI(net233));
 sg13g2_tiehi _5005__234 (.L_HI(net234));
 sg13g2_tiehi _5004__235 (.L_HI(net235));
 sg13g2_tiehi _5113__236 (.L_HI(net236));
 sg13g2_tiehi _5003__237 (.L_HI(net237));
 sg13g2_tiehi _5161__238 (.L_HI(net238));
 sg13g2_tiehi _5002__239 (.L_HI(net239));
 sg13g2_tiehi _5112__240 (.L_HI(net240));
 sg13g2_tiehi _5001__241 (.L_HI(net241));
 sg13g2_tiehi _5185__242 (.L_HI(net242));
 sg13g2_tiehi _5000__243 (.L_HI(net243));
 sg13g2_tiehi _5111__244 (.L_HI(net244));
 sg13g2_tiehi _4999__245 (.L_HI(net245));
 sg13g2_tiehi _5160__246 (.L_HI(net246));
 sg13g2_tiehi _4998__247 (.L_HI(net247));
 sg13g2_tiehi _5110__248 (.L_HI(net248));
 sg13g2_tiehi _4997__249 (.L_HI(net249));
 sg13g2_tiehi _5206__250 (.L_HI(net250));
 sg13g2_tiehi _4996__251 (.L_HI(net251));
 sg13g2_tiehi _5109__252 (.L_HI(net252));
 sg13g2_tiehi _4995__253 (.L_HI(net253));
 sg13g2_tiehi _5159__254 (.L_HI(net254));
 sg13g2_tiehi _4994__255 (.L_HI(net255));
 sg13g2_tiehi _5108__256 (.L_HI(net256));
 sg13g2_tiehi _4993__257 (.L_HI(net257));
 sg13g2_tiehi _5184__258 (.L_HI(net258));
 sg13g2_tiehi _4992__259 (.L_HI(net259));
 sg13g2_tiehi _5107__260 (.L_HI(net260));
 sg13g2_tiehi _4834__261 (.L_HI(net261));
 sg13g2_tiehi _5064__262 (.L_HI(net262));
 sg13g2_tiehi _5065__263 (.L_HI(net263));
 sg13g2_tiehi _5066__264 (.L_HI(net264));
 sg13g2_tiehi _4991__265 (.L_HI(net265));
 sg13g2_tiehi _5158__266 (.L_HI(net266));
 sg13g2_tiehi _4990__267 (.L_HI(net267));
 sg13g2_tiehi _5106__268 (.L_HI(net268));
 sg13g2_tiehi _4989__269 (.L_HI(net269));
 sg13g2_tiehi _4988__270 (.L_HI(net270));
 sg13g2_tiehi _5105__271 (.L_HI(net271));
 sg13g2_tiehi _4987__272 (.L_HI(net272));
 sg13g2_tiehi _5157__273 (.L_HI(net273));
 sg13g2_tiehi _4986__274 (.L_HI(net274));
 sg13g2_tiehi _5104__275 (.L_HI(net275));
 sg13g2_tiehi _4985__276 (.L_HI(net276));
 sg13g2_tiehi _5183__277 (.L_HI(net277));
 sg13g2_tiehi _4984__278 (.L_HI(net278));
 sg13g2_tiehi _5103__279 (.L_HI(net279));
 sg13g2_tiehi _4983__280 (.L_HI(net280));
 sg13g2_tiehi _5156__281 (.L_HI(net281));
 sg13g2_tiehi _4982__282 (.L_HI(net282));
 sg13g2_tiehi _5102__283 (.L_HI(net283));
 sg13g2_tiehi _4981__284 (.L_HI(net284));
 sg13g2_tiehi _5205__285 (.L_HI(net285));
 sg13g2_tiehi _4980__286 (.L_HI(net286));
 sg13g2_tiehi _5101__287 (.L_HI(net287));
 sg13g2_tiehi _4979__288 (.L_HI(net288));
 sg13g2_tiehi _5155__289 (.L_HI(net289));
 sg13g2_tiehi _4978__290 (.L_HI(net290));
 sg13g2_tiehi _5100__291 (.L_HI(net291));
 sg13g2_tiehi _4977__292 (.L_HI(net292));
 sg13g2_tiehi _5182__293 (.L_HI(net293));
 sg13g2_tiehi _4976__294 (.L_HI(net294));
 sg13g2_tiehi _5099__295 (.L_HI(net295));
 sg13g2_tiehi _4975__296 (.L_HI(net296));
 sg13g2_tiehi _5154__297 (.L_HI(net297));
 sg13g2_tiehi _4974__298 (.L_HI(net298));
 sg13g2_tiehi _5098__299 (.L_HI(net299));
 sg13g2_tiehi _4973__300 (.L_HI(net300));
 sg13g2_tiehi _4972__301 (.L_HI(net301));
 sg13g2_tiehi _5097__302 (.L_HI(net302));
 sg13g2_tiehi _4971__303 (.L_HI(net303));
 sg13g2_tiehi _5153__304 (.L_HI(net304));
 sg13g2_tiehi _4970__305 (.L_HI(net305));
 sg13g2_tiehi _5096__306 (.L_HI(net306));
 sg13g2_tiehi _4969__307 (.L_HI(net307));
 sg13g2_tiehi _5181__308 (.L_HI(net308));
 sg13g2_tiehi _4968__309 (.L_HI(net309));
 sg13g2_tiehi _5095__310 (.L_HI(net310));
 sg13g2_tiehi _4967__311 (.L_HI(net311));
 sg13g2_tiehi _5152__312 (.L_HI(net312));
 sg13g2_tiehi _4966__313 (.L_HI(net313));
 sg13g2_tiehi _5094__314 (.L_HI(net314));
 sg13g2_tiehi _4965__315 (.L_HI(net315));
 sg13g2_tiehi _5204__316 (.L_HI(net316));
 sg13g2_tiehi _4964__317 (.L_HI(net317));
 sg13g2_tiehi _5093__318 (.L_HI(net318));
 sg13g2_tiehi _4963__319 (.L_HI(net319));
 sg13g2_tiehi _5151__320 (.L_HI(net320));
 sg13g2_tiehi _4962__321 (.L_HI(net321));
 sg13g2_tiehi _5092__322 (.L_HI(net322));
 sg13g2_tiehi _4961__323 (.L_HI(net323));
 sg13g2_tiehi _4960__324 (.L_HI(net324));
 sg13g2_tiehi _4959__325 (.L_HI(net325));
 sg13g2_tiehi _4958__326 (.L_HI(net326));
 sg13g2_tiehi _4957__327 (.L_HI(net327));
 sg13g2_tiehi _4956__328 (.L_HI(net328));
 sg13g2_tiehi _4955__329 (.L_HI(net329));
 sg13g2_tiehi _4954__330 (.L_HI(net330));
 sg13g2_tiehi _4953__331 (.L_HI(net331));
 sg13g2_tiehi _4952__332 (.L_HI(net332));
 sg13g2_tiehi _4951__333 (.L_HI(net333));
 sg13g2_tiehi _4950__334 (.L_HI(net334));
 sg13g2_tiehi _4949__335 (.L_HI(net335));
 sg13g2_tiehi _4948__336 (.L_HI(net336));
 sg13g2_tiehi _4947__337 (.L_HI(net337));
 sg13g2_tiehi _4946__338 (.L_HI(net338));
 sg13g2_tiehi _4945__339 (.L_HI(net339));
 sg13g2_tiehi _4944__340 (.L_HI(net340));
 sg13g2_tiehi _4943__341 (.L_HI(net341));
 sg13g2_tiehi _4942__342 (.L_HI(net342));
 sg13g2_tiehi _4941__343 (.L_HI(net343));
 sg13g2_tiehi _4940__344 (.L_HI(net344));
 sg13g2_tiehi _4939__345 (.L_HI(net345));
 sg13g2_tiehi _4938__346 (.L_HI(net346));
 sg13g2_tiehi _5180__347 (.L_HI(net347));
 sg13g2_tiehi _4937__348 (.L_HI(net348));
 sg13g2_tiehi _5091__349 (.L_HI(net349));
 sg13g2_tiehi _4936__350 (.L_HI(net350));
 sg13g2_tiehi _5150__351 (.L_HI(net351));
 sg13g2_tiehi _4935__352 (.L_HI(net352));
 sg13g2_tiehi _5090__353 (.L_HI(net353));
 sg13g2_tiehi _4934__354 (.L_HI(net354));
 sg13g2_tiehi _5089__355 (.L_HI(net355));
 sg13g2_tiehi _4933__356 (.L_HI(net356));
 sg13g2_tiehi _5088__357 (.L_HI(net357));
 sg13g2_tiehi _4932__358 (.L_HI(net358));
 sg13g2_tiehi _5087__359 (.L_HI(net359));
 sg13g2_tiehi _4931__360 (.L_HI(net360));
 sg13g2_tiehi _5086__361 (.L_HI(net361));
 sg13g2_tiehi _4930__362 (.L_HI(net362));
 sg13g2_tiehi _5085__363 (.L_HI(net363));
 sg13g2_tiehi _4929__364 (.L_HI(net364));
 sg13g2_tiehi _5084__365 (.L_HI(net365));
 sg13g2_tiehi _4928__366 (.L_HI(net366));
 sg13g2_tiehi _5083__367 (.L_HI(net367));
 sg13g2_tiehi _4927__368 (.L_HI(net368));
 sg13g2_tiehi _5082__369 (.L_HI(net369));
 sg13g2_tiehi _4926__370 (.L_HI(net370));
 sg13g2_tiehi _5081__371 (.L_HI(net371));
 sg13g2_tiehi _4925__372 (.L_HI(net372));
 sg13g2_tiehi _5203__373 (.L_HI(net373));
 sg13g2_tiehi _4924__374 (.L_HI(net374));
 sg13g2_tiehi _5080__375 (.L_HI(net375));
 sg13g2_tiehi _4923__376 (.L_HI(net376));
 sg13g2_tiehi _5149__377 (.L_HI(net377));
 sg13g2_tiehi _4922__378 (.L_HI(net378));
 sg13g2_tiehi _5079__379 (.L_HI(net379));
 sg13g2_tiehi _4921__380 (.L_HI(net380));
 sg13g2_tiehi _5179__381 (.L_HI(net381));
 sg13g2_tiehi _4920__382 (.L_HI(net382));
 sg13g2_tiehi _5078__383 (.L_HI(net383));
 sg13g2_tiehi _4919__384 (.L_HI(net384));
 sg13g2_tiehi _5148__385 (.L_HI(net385));
 sg13g2_tiehi _4918__386 (.L_HI(net386));
 sg13g2_tiehi _5077__387 (.L_HI(net387));
 sg13g2_tiehi _4917__388 (.L_HI(net388));
 sg13g2_tiehi _5202__389 (.L_HI(net389));
 sg13g2_tiehi _4916__390 (.L_HI(net390));
 sg13g2_tiehi _5076__391 (.L_HI(net391));
 sg13g2_tiehi _4915__392 (.L_HI(net392));
 sg13g2_tiehi _5147__393 (.L_HI(net393));
 sg13g2_tiehi _4914__394 (.L_HI(net394));
 sg13g2_tiehi _5075__395 (.L_HI(net395));
 sg13g2_tiehi _4913__396 (.L_HI(net396));
 sg13g2_tiehi _5178__397 (.L_HI(net397));
 sg13g2_tiehi _4912__398 (.L_HI(net398));
 sg13g2_tiehi _5074__399 (.L_HI(net399));
 sg13g2_tiehi _4911__400 (.L_HI(net400));
 sg13g2_tiehi _5146__401 (.L_HI(net401));
 sg13g2_tiehi _5067__402 (.L_HI(net402));
 sg13g2_tiehi _5207__403 (.L_HI(net403));
 sg13g2_tiehi _4910__404 (.L_HI(net404));
 sg13g2_inv_1 _2612__1 (.Y(net405),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo heichips25_bagel_20 (.L_LO(net20));
 sg13g2_tielo heichips25_bagel_21 (.L_LO(net21));
 sg13g2_tielo heichips25_bagel_22 (.L_LO(net22));
 sg13g2_tielo heichips25_bagel_23 (.L_LO(net23));
 sg13g2_tielo heichips25_bagel_24 (.L_LO(net24));
 sg13g2_tielo heichips25_bagel_25 (.L_LO(net25));
 sg13g2_tielo heichips25_bagel_26 (.L_LO(net26));
 sg13g2_tielo heichips25_bagel_27 (.L_LO(net27));
 sg13g2_tielo heichips25_bagel_28 (.L_LO(net28));
 sg13g2_tielo heichips25_bagel_29 (.L_LO(net29));
 sg13g2_tielo heichips25_bagel_30 (.L_LO(net30));
 sg13g2_tiehi _5073__31 (.L_HI(net31));
 sg13g2_buf_8 fanout544 (.A(_1089_),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(_0691_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_0691_),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(_0881_),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(_0881_),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(_0682_),
    .X(net549));
 sg13g2_buf_8 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_1 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_1 fanout552 (.A(net555),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_8 fanout555 (.A(_1300_),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(net560),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(net560),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(net560),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_8 fanout560 (.A(_1300_),
    .X(net560));
 sg13g2_buf_8 fanout561 (.A(net565),
    .X(net561));
 sg13g2_buf_1 fanout562 (.A(net565),
    .X(net562));
 sg13g2_buf_8 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(_1303_),
    .X(net565));
 sg13g2_buf_8 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(net570),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(net570),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(_1303_),
    .X(net570));
 sg13g2_buf_8 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(_0853_),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(net577),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(net577),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(_0702_),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(net582),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net582),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(_0702_),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_0701_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_8 fanout585 (.A(net587),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(_0687_),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(net592),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net592),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(net592),
    .X(net590));
 sg13g2_buf_1 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(_0687_),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(_0686_),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(_0659_),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(_0645_),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(_0645_),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(_0645_),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(\tmds_green.n132 ),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(\tmds_green.n100 ),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(\tmds_blue.n100 ),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(net607),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(display_enable),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(\videogen.fancy_shader.video_y[0] ),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(\videogen.fancy_shader.n646[8] ),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[5] ),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(net613),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[4] ),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[3] ),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(net620),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(net627),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(net627),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(net627),
    .X(net625));
 sg13g2_buf_1 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[2] ),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(\videogen.test_lut_thingy.pixel_feeder_inst.h_pix[0] ),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(\videogen.fancy_shader.video_x[7] ),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net648),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net640),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net640),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(net640),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net640),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net640),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_1 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net648),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net643),
    .X(net641));
 sg13g2_buf_1 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net646),
    .X(net643));
 sg13g2_buf_8 fanout644 (.A(net646),
    .X(net644));
 sg13g2_buf_1 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_8 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(clk_video),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net651),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net654),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_1 fanout654 (.A(net672),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net659),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(net659),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net672),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(net662),
    .X(net660));
 sg13g2_buf_1 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(net672),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net666),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net666),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(net672),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net671),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net671),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_8 fanout672 (.A(net693),
    .X(net672));
 sg13g2_buf_8 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net682),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(net682),
    .X(net675));
 sg13g2_buf_1 fanout676 (.A(net682),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net682),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(net682),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net681),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net693),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(net687),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net693),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(net692),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net692),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(\clockdiv.q2temp ),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(net700),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net699),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(net699),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net446),
    .X(net700));
 sg13g2_buf_8 fanout701 (.A(net703),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(net706),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(net724),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(net711),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(net711),
    .X(net709));
 sg13g2_buf_1 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net724),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(net714),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(net724),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(net718),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(net718),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(net724),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net723),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(net723),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net744),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net733),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net733),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net733),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(net732),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net732),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net744),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net738),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net738),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net744),
    .X(net738));
 sg13g2_buf_8 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(net743),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(\clockdiv.q1 ),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(net751),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_8 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(_0658_),
    .X(net751));
 sg13g2_buf_8 fanout752 (.A(net756),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net756),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(ui_in[7]),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net761),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net761),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(net761),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(ui_in[7]),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net766),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net766),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net766),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net772),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(net769),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net772),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_8 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(ui_in[6]),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(ui_in[5]),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net778),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(net778),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(ui_in[5]),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net783),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net783),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net783),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(ui_in[5]),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net794),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net788),
    .X(net786));
 sg13g2_buf_1 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net794),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net793),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(ui_in[4]),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(rst_n),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net806),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net806),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(net806),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(net805),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(net805),
    .X(net804));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(rst_n),
    .X(net806));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(tmds_b));
 sg13g2_buf_1 output4 (.A(net4),
    .X(tmds_clk));
 sg13g2_buf_1 output5 (.A(net5),
    .X(tmds_g));
 sg13g2_buf_1 output6 (.A(net6),
    .X(tmds_r));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_bagel_19 (.L_LO(net19));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\clockdiv.q2 ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0623_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold3 (.A(\serialize.n420[2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold4 (.A(\serialize.n420[3] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold5 (.A(\serialize.n420[0] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold6 (.A(\serialize.n420[1] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold7 (.A(\serialize.bit_cnt[0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold8 (.A(\serialize.n420[4] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold9 (.A(\serialize.n414[1] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0004_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0262_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold12 (.A(\serialize.n414[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold13 (.A(\serialize.n414[5] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold14 (.A(\serialize.n420[6] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold15 (.A(\serialize.n431[6] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold16 (.A(\serialize.n411[0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold17 (.A(\serialize.n411[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold18 (.A(\serialize.n414[0] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold19 (.A(\serialize.n411[3] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold20 (.A(\serialize.n417[7] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold21 (.A(\serialize.n411[5] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold22 (.A(\serialize.n417[5] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold23 (.A(\serialize.n417[0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold24 (.A(\serialize.n414[6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold25 (.A(\serialize.n411[6] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold26 (.A(\serialize.n411[7] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold27 (.A(\clockdiv.q0 ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold28 (.A(\serialize.n417[3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold29 (.A(\serialize.n429[3] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold30 (.A(\serialize.n417[6] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold31 (.A(\serialize.n414[2] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold32 (.A(\serialize.n417[2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold33 (.A(\serialize.n414[7] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold34 (.A(\serialize.n414[4] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold35 (.A(\serialize.n417[1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold36 (.A(\serialize.n411[1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold37 (.A(\serialize.n411[4] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold38 (.A(\serialize.n417[4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold39 (.A(\serialize.n429[4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold40 (.A(\serialize.bit_cnt[1] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold41 (.A(\serialize.n410 ),
    .X(net446));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_41 ();
 sg13g2_fill_2 FILLER_0_48 ();
 sg13g2_fill_1 FILLER_0_55 ();
 sg13g2_decap_8 FILLER_0_60 ();
 sg13g2_decap_8 FILLER_0_67 ();
 sg13g2_fill_1 FILLER_0_74 ();
 sg13g2_decap_4 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_94 ();
 sg13g2_decap_4 FILLER_0_101 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_4 FILLER_0_126 ();
 sg13g2_decap_4 FILLER_0_135 ();
 sg13g2_fill_2 FILLER_0_139 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_4 FILLER_0_179 ();
 sg13g2_fill_2 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_4 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_fill_2 FILLER_0_227 ();
 sg13g2_fill_1 FILLER_0_229 ();
 sg13g2_fill_1 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_317 ();
 sg13g2_fill_2 FILLER_0_328 ();
 sg13g2_decap_4 FILLER_0_334 ();
 sg13g2_fill_1 FILLER_0_338 ();
 sg13g2_decap_4 FILLER_0_349 ();
 sg13g2_fill_1 FILLER_0_353 ();
 sg13g2_decap_4 FILLER_0_358 ();
 sg13g2_fill_1 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_fill_2 FILLER_0_408 ();
 sg13g2_fill_1 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_decap_8 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_decap_8 FILLER_0_453 ();
 sg13g2_decap_8 FILLER_0_460 ();
 sg13g2_decap_8 FILLER_0_467 ();
 sg13g2_decap_8 FILLER_0_474 ();
 sg13g2_decap_8 FILLER_0_494 ();
 sg13g2_decap_8 FILLER_0_501 ();
 sg13g2_decap_8 FILLER_0_508 ();
 sg13g2_decap_8 FILLER_0_515 ();
 sg13g2_decap_8 FILLER_0_522 ();
 sg13g2_decap_8 FILLER_0_529 ();
 sg13g2_decap_8 FILLER_0_536 ();
 sg13g2_decap_8 FILLER_0_543 ();
 sg13g2_decap_8 FILLER_0_550 ();
 sg13g2_decap_8 FILLER_0_557 ();
 sg13g2_decap_8 FILLER_0_564 ();
 sg13g2_decap_8 FILLER_0_571 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_4 FILLER_0_616 ();
 sg13g2_fill_1 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_641 ();
 sg13g2_decap_8 FILLER_0_648 ();
 sg13g2_decap_4 FILLER_0_655 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_8 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_decap_8 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_8 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_decap_8 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_fill_2 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_65 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_fill_1 FILLER_1_195 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_313 ();
 sg13g2_fill_1 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_370 ();
 sg13g2_decap_4 FILLER_1_425 ();
 sg13g2_decap_8 FILLER_1_508 ();
 sg13g2_decap_8 FILLER_1_515 ();
 sg13g2_decap_8 FILLER_1_522 ();
 sg13g2_decap_8 FILLER_1_529 ();
 sg13g2_decap_8 FILLER_1_536 ();
 sg13g2_decap_8 FILLER_1_543 ();
 sg13g2_decap_8 FILLER_1_550 ();
 sg13g2_decap_8 FILLER_1_557 ();
 sg13g2_decap_8 FILLER_1_564 ();
 sg13g2_fill_2 FILLER_1_571 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_fill_1 FILLER_1_611 ();
 sg13g2_fill_1 FILLER_1_629 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_fill_1 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_decap_8 FILLER_1_731 ();
 sg13g2_decap_8 FILLER_1_738 ();
 sg13g2_fill_2 FILLER_1_745 ();
 sg13g2_fill_1 FILLER_1_747 ();
 sg13g2_decap_8 FILLER_1_753 ();
 sg13g2_decap_8 FILLER_1_760 ();
 sg13g2_decap_8 FILLER_1_767 ();
 sg13g2_decap_8 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_879 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_decap_8 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_942 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_977 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_decap_8 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_fill_2 FILLER_1_1026 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_4 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_66 ();
 sg13g2_fill_2 FILLER_2_73 ();
 sg13g2_fill_1 FILLER_2_75 ();
 sg13g2_decap_8 FILLER_2_99 ();
 sg13g2_decap_8 FILLER_2_106 ();
 sg13g2_decap_4 FILLER_2_113 ();
 sg13g2_fill_2 FILLER_2_117 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_4 FILLER_2_134 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_decap_8 FILLER_2_209 ();
 sg13g2_decap_4 FILLER_2_216 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_decap_4 FILLER_2_231 ();
 sg13g2_fill_2 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_fill_1 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_278 ();
 sg13g2_fill_2 FILLER_2_285 ();
 sg13g2_fill_1 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_309 ();
 sg13g2_decap_4 FILLER_2_316 ();
 sg13g2_fill_1 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_4 FILLER_2_343 ();
 sg13g2_fill_1 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_4 FILLER_2_441 ();
 sg13g2_decap_4 FILLER_2_472 ();
 sg13g2_decap_8 FILLER_2_519 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_4 FILLER_2_574 ();
 sg13g2_fill_2 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_597 ();
 sg13g2_fill_1 FILLER_2_604 ();
 sg13g2_decap_8 FILLER_2_614 ();
 sg13g2_fill_2 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_643 ();
 sg13g2_fill_1 FILLER_2_650 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_4 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_684 ();
 sg13g2_fill_2 FILLER_2_691 ();
 sg13g2_decap_4 FILLER_2_701 ();
 sg13g2_fill_2 FILLER_2_710 ();
 sg13g2_decap_4 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_761 ();
 sg13g2_decap_8 FILLER_2_768 ();
 sg13g2_decap_8 FILLER_2_775 ();
 sg13g2_decap_8 FILLER_2_782 ();
 sg13g2_decap_8 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_803 ();
 sg13g2_decap_8 FILLER_2_810 ();
 sg13g2_decap_8 FILLER_2_817 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_decap_8 FILLER_2_859 ();
 sg13g2_decap_8 FILLER_2_866 ();
 sg13g2_decap_8 FILLER_2_873 ();
 sg13g2_decap_8 FILLER_2_880 ();
 sg13g2_decap_8 FILLER_2_887 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_decap_8 FILLER_2_985 ();
 sg13g2_decap_8 FILLER_2_992 ();
 sg13g2_decap_8 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1013 ();
 sg13g2_decap_8 FILLER_2_1020 ();
 sg13g2_fill_2 FILLER_2_1027 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_26 ();
 sg13g2_fill_1 FILLER_3_33 ();
 sg13g2_decap_4 FILLER_3_38 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_58 ();
 sg13g2_decap_8 FILLER_3_65 ();
 sg13g2_fill_2 FILLER_3_72 ();
 sg13g2_fill_1 FILLER_3_74 ();
 sg13g2_fill_1 FILLER_3_85 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_98 ();
 sg13g2_fill_1 FILLER_3_100 ();
 sg13g2_decap_8 FILLER_3_118 ();
 sg13g2_decap_8 FILLER_3_125 ();
 sg13g2_decap_8 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_166 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_fill_2 FILLER_3_180 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_4 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_fill_1 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_346 ();
 sg13g2_decap_4 FILLER_3_351 ();
 sg13g2_fill_2 FILLER_3_372 ();
 sg13g2_fill_2 FILLER_3_405 ();
 sg13g2_decap_4 FILLER_3_444 ();
 sg13g2_fill_2 FILLER_3_461 ();
 sg13g2_fill_1 FILLER_3_463 ();
 sg13g2_decap_8 FILLER_3_468 ();
 sg13g2_decap_8 FILLER_3_475 ();
 sg13g2_decap_4 FILLER_3_492 ();
 sg13g2_fill_1 FILLER_3_496 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_fill_1 FILLER_3_515 ();
 sg13g2_fill_1 FILLER_3_521 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_fill_1 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_555 ();
 sg13g2_decap_8 FILLER_3_562 ();
 sg13g2_decap_8 FILLER_3_569 ();
 sg13g2_decap_8 FILLER_3_576 ();
 sg13g2_decap_4 FILLER_3_583 ();
 sg13g2_decap_4 FILLER_3_591 ();
 sg13g2_fill_1 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_fill_2 FILLER_3_644 ();
 sg13g2_fill_1 FILLER_3_674 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_decap_4 FILLER_3_698 ();
 sg13g2_fill_2 FILLER_3_715 ();
 sg13g2_fill_1 FILLER_3_717 ();
 sg13g2_fill_2 FILLER_3_733 ();
 sg13g2_fill_1 FILLER_3_735 ();
 sg13g2_fill_2 FILLER_3_771 ();
 sg13g2_fill_1 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_8 FILLER_3_913 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_decap_8 FILLER_3_927 ();
 sg13g2_decap_8 FILLER_3_934 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_8 FILLER_3_976 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_4_8 ();
 sg13g2_fill_2 FILLER_4_15 ();
 sg13g2_decap_8 FILLER_4_45 ();
 sg13g2_decap_8 FILLER_4_52 ();
 sg13g2_decap_4 FILLER_4_59 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_69 ();
 sg13g2_decap_4 FILLER_4_76 ();
 sg13g2_fill_2 FILLER_4_80 ();
 sg13g2_decap_4 FILLER_4_86 ();
 sg13g2_fill_2 FILLER_4_90 ();
 sg13g2_fill_2 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_149 ();
 sg13g2_decap_4 FILLER_4_156 ();
 sg13g2_decap_4 FILLER_4_183 ();
 sg13g2_fill_1 FILLER_4_187 ();
 sg13g2_decap_4 FILLER_4_192 ();
 sg13g2_fill_1 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_201 ();
 sg13g2_decap_8 FILLER_4_208 ();
 sg13g2_decap_4 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_219 ();
 sg13g2_fill_2 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_fill_1 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_fill_2 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_fill_2 FILLER_4_459 ();
 sg13g2_fill_1 FILLER_4_461 ();
 sg13g2_decap_8 FILLER_4_489 ();
 sg13g2_decap_8 FILLER_4_496 ();
 sg13g2_decap_8 FILLER_4_503 ();
 sg13g2_decap_4 FILLER_4_510 ();
 sg13g2_fill_2 FILLER_4_514 ();
 sg13g2_fill_2 FILLER_4_543 ();
 sg13g2_fill_1 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_614 ();
 sg13g2_decap_8 FILLER_4_621 ();
 sg13g2_decap_8 FILLER_4_628 ();
 sg13g2_fill_1 FILLER_4_635 ();
 sg13g2_decap_8 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_652 ();
 sg13g2_decap_4 FILLER_4_659 ();
 sg13g2_fill_1 FILLER_4_663 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_fill_2 FILLER_4_700 ();
 sg13g2_fill_1 FILLER_4_702 ();
 sg13g2_decap_4 FILLER_4_708 ();
 sg13g2_fill_2 FILLER_4_712 ();
 sg13g2_fill_1 FILLER_4_719 ();
 sg13g2_decap_8 FILLER_4_730 ();
 sg13g2_decap_8 FILLER_4_737 ();
 sg13g2_fill_1 FILLER_4_744 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_4 FILLER_4_768 ();
 sg13g2_decap_8 FILLER_4_794 ();
 sg13g2_decap_4 FILLER_4_801 ();
 sg13g2_fill_1 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_8 FILLER_4_834 ();
 sg13g2_decap_8 FILLER_4_841 ();
 sg13g2_decap_8 FILLER_4_848 ();
 sg13g2_decap_8 FILLER_4_855 ();
 sg13g2_decap_8 FILLER_4_862 ();
 sg13g2_decap_8 FILLER_4_869 ();
 sg13g2_decap_8 FILLER_4_876 ();
 sg13g2_decap_8 FILLER_4_883 ();
 sg13g2_decap_8 FILLER_4_890 ();
 sg13g2_decap_8 FILLER_4_897 ();
 sg13g2_decap_8 FILLER_4_904 ();
 sg13g2_decap_8 FILLER_4_911 ();
 sg13g2_decap_8 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_925 ();
 sg13g2_decap_8 FILLER_4_932 ();
 sg13g2_decap_8 FILLER_4_939 ();
 sg13g2_decap_8 FILLER_4_946 ();
 sg13g2_decap_8 FILLER_4_953 ();
 sg13g2_decap_8 FILLER_4_960 ();
 sg13g2_decap_8 FILLER_4_967 ();
 sg13g2_decap_8 FILLER_4_974 ();
 sg13g2_decap_8 FILLER_4_981 ();
 sg13g2_decap_8 FILLER_4_988 ();
 sg13g2_decap_8 FILLER_4_995 ();
 sg13g2_decap_8 FILLER_4_1002 ();
 sg13g2_decap_8 FILLER_4_1009 ();
 sg13g2_decap_8 FILLER_4_1016 ();
 sg13g2_decap_4 FILLER_4_1023 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_decap_8 FILLER_5_30 ();
 sg13g2_decap_8 FILLER_5_37 ();
 sg13g2_decap_8 FILLER_5_44 ();
 sg13g2_decap_4 FILLER_5_51 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_fill_2 FILLER_5_104 ();
 sg13g2_fill_1 FILLER_5_106 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_150 ();
 sg13g2_fill_2 FILLER_5_173 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_4 FILLER_5_299 ();
 sg13g2_fill_2 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_309 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_decap_4 FILLER_5_334 ();
 sg13g2_fill_2 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_decap_4 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_5_465 ();
 sg13g2_decap_4 FILLER_5_471 ();
 sg13g2_fill_2 FILLER_5_479 ();
 sg13g2_fill_1 FILLER_5_481 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_fill_2 FILLER_5_504 ();
 sg13g2_fill_1 FILLER_5_506 ();
 sg13g2_fill_2 FILLER_5_541 ();
 sg13g2_fill_1 FILLER_5_543 ();
 sg13g2_fill_2 FILLER_5_549 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_fill_1 FILLER_5_585 ();
 sg13g2_fill_2 FILLER_5_599 ();
 sg13g2_decap_4 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_614 ();
 sg13g2_decap_4 FILLER_5_621 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_659 ();
 sg13g2_fill_2 FILLER_5_666 ();
 sg13g2_fill_2 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_fill_1 FILLER_5_686 ();
 sg13g2_fill_2 FILLER_5_713 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_fill_2 FILLER_5_746 ();
 sg13g2_decap_4 FILLER_5_753 ();
 sg13g2_fill_2 FILLER_5_757 ();
 sg13g2_decap_8 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_fill_1 FILLER_5_778 ();
 sg13g2_fill_2 FILLER_5_785 ();
 sg13g2_decap_4 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_4 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_4 FILLER_6_4 ();
 sg13g2_fill_1 FILLER_6_8 ();
 sg13g2_fill_2 FILLER_6_13 ();
 sg13g2_fill_1 FILLER_6_15 ();
 sg13g2_decap_8 FILLER_6_24 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_fill_2 FILLER_6_135 ();
 sg13g2_fill_2 FILLER_6_170 ();
 sg13g2_decap_4 FILLER_6_176 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_202 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_fill_2 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_268 ();
 sg13g2_fill_2 FILLER_6_327 ();
 sg13g2_fill_2 FILLER_6_335 ();
 sg13g2_fill_1 FILLER_6_337 ();
 sg13g2_fill_2 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_fill_2 FILLER_6_388 ();
 sg13g2_fill_1 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_401 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_1 FILLER_6_409 ();
 sg13g2_decap_4 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_6_430 ();
 sg13g2_decap_4 FILLER_6_437 ();
 sg13g2_fill_2 FILLER_6_441 ();
 sg13g2_fill_1 FILLER_6_470 ();
 sg13g2_decap_4 FILLER_6_508 ();
 sg13g2_decap_4 FILLER_6_520 ();
 sg13g2_fill_2 FILLER_6_524 ();
 sg13g2_decap_4 FILLER_6_562 ();
 sg13g2_fill_2 FILLER_6_594 ();
 sg13g2_decap_4 FILLER_6_600 ();
 sg13g2_decap_8 FILLER_6_611 ();
 sg13g2_decap_8 FILLER_6_618 ();
 sg13g2_decap_4 FILLER_6_625 ();
 sg13g2_fill_1 FILLER_6_629 ();
 sg13g2_fill_2 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_644 ();
 sg13g2_decap_4 FILLER_6_658 ();
 sg13g2_fill_1 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_677 ();
 sg13g2_decap_4 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_688 ();
 sg13g2_decap_4 FILLER_6_697 ();
 sg13g2_decap_4 FILLER_6_706 ();
 sg13g2_fill_2 FILLER_6_710 ();
 sg13g2_decap_4 FILLER_6_722 ();
 sg13g2_fill_1 FILLER_6_732 ();
 sg13g2_decap_4 FILLER_6_737 ();
 sg13g2_fill_2 FILLER_6_769 ();
 sg13g2_fill_1 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_fill_2 FILLER_6_803 ();
 sg13g2_fill_1 FILLER_6_805 ();
 sg13g2_fill_1 FILLER_6_814 ();
 sg13g2_fill_1 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_843 ();
 sg13g2_fill_2 FILLER_6_850 ();
 sg13g2_fill_1 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_872 ();
 sg13g2_decap_8 FILLER_6_879 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_4 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_51 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_2 FILLER_7_62 ();
 sg13g2_decap_8 FILLER_7_68 ();
 sg13g2_decap_8 FILLER_7_75 ();
 sg13g2_decap_8 FILLER_7_82 ();
 sg13g2_decap_8 FILLER_7_89 ();
 sg13g2_decap_8 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_103 ();
 sg13g2_fill_1 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_114 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_142 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_4 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_decap_4 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_289 ();
 sg13g2_decap_8 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_decap_4 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_4 FILLER_7_352 ();
 sg13g2_fill_2 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_fill_1 FILLER_7_386 ();
 sg13g2_decap_4 FILLER_7_439 ();
 sg13g2_decap_8 FILLER_7_464 ();
 sg13g2_fill_2 FILLER_7_471 ();
 sg13g2_decap_8 FILLER_7_477 ();
 sg13g2_fill_2 FILLER_7_484 ();
 sg13g2_decap_8 FILLER_7_496 ();
 sg13g2_decap_8 FILLER_7_503 ();
 sg13g2_decap_4 FILLER_7_510 ();
 sg13g2_fill_2 FILLER_7_514 ();
 sg13g2_decap_8 FILLER_7_522 ();
 sg13g2_fill_2 FILLER_7_529 ();
 sg13g2_decap_4 FILLER_7_536 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_565 ();
 sg13g2_fill_1 FILLER_7_576 ();
 sg13g2_fill_1 FILLER_7_590 ();
 sg13g2_fill_1 FILLER_7_601 ();
 sg13g2_fill_1 FILLER_7_619 ();
 sg13g2_fill_2 FILLER_7_633 ();
 sg13g2_fill_1 FILLER_7_635 ();
 sg13g2_fill_2 FILLER_7_668 ();
 sg13g2_decap_4 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_fill_2 FILLER_7_721 ();
 sg13g2_fill_2 FILLER_7_753 ();
 sg13g2_fill_1 FILLER_7_755 ();
 sg13g2_fill_2 FILLER_7_768 ();
 sg13g2_fill_1 FILLER_7_770 ();
 sg13g2_fill_2 FILLER_7_775 ();
 sg13g2_fill_1 FILLER_7_781 ();
 sg13g2_decap_4 FILLER_7_787 ();
 sg13g2_decap_8 FILLER_7_799 ();
 sg13g2_decap_4 FILLER_7_806 ();
 sg13g2_fill_1 FILLER_7_810 ();
 sg13g2_decap_4 FILLER_7_842 ();
 sg13g2_fill_1 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_878 ();
 sg13g2_decap_8 FILLER_7_885 ();
 sg13g2_decap_8 FILLER_7_892 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_906 ();
 sg13g2_decap_8 FILLER_7_913 ();
 sg13g2_decap_8 FILLER_7_920 ();
 sg13g2_decap_8 FILLER_7_927 ();
 sg13g2_decap_8 FILLER_7_934 ();
 sg13g2_decap_8 FILLER_7_941 ();
 sg13g2_decap_8 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_955 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_decap_8 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1004 ();
 sg13g2_decap_8 FILLER_7_1011 ();
 sg13g2_decap_8 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_decap_8 FILLER_8_20 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_fill_1 FILLER_8_81 ();
 sg13g2_fill_2 FILLER_8_92 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_142 ();
 sg13g2_fill_1 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_150 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_194 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_4 FILLER_8_237 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_decap_4 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_257 ();
 sg13g2_decap_4 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_292 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_4 FILLER_8_349 ();
 sg13g2_fill_2 FILLER_8_362 ();
 sg13g2_fill_1 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_fill_2 FILLER_8_376 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_411 ();
 sg13g2_decap_4 FILLER_8_418 ();
 sg13g2_fill_2 FILLER_8_422 ();
 sg13g2_decap_8 FILLER_8_433 ();
 sg13g2_decap_8 FILLER_8_440 ();
 sg13g2_decap_4 FILLER_8_447 ();
 sg13g2_fill_1 FILLER_8_451 ();
 sg13g2_fill_2 FILLER_8_474 ();
 sg13g2_decap_8 FILLER_8_520 ();
 sg13g2_decap_8 FILLER_8_527 ();
 sg13g2_decap_8 FILLER_8_534 ();
 sg13g2_fill_2 FILLER_8_541 ();
 sg13g2_fill_1 FILLER_8_543 ();
 sg13g2_fill_1 FILLER_8_579 ();
 sg13g2_decap_8 FILLER_8_593 ();
 sg13g2_fill_2 FILLER_8_600 ();
 sg13g2_fill_1 FILLER_8_602 ();
 sg13g2_fill_2 FILLER_8_608 ();
 sg13g2_fill_1 FILLER_8_610 ();
 sg13g2_decap_8 FILLER_8_626 ();
 sg13g2_fill_2 FILLER_8_633 ();
 sg13g2_fill_1 FILLER_8_635 ();
 sg13g2_fill_1 FILLER_8_640 ();
 sg13g2_decap_4 FILLER_8_645 ();
 sg13g2_decap_8 FILLER_8_654 ();
 sg13g2_decap_8 FILLER_8_661 ();
 sg13g2_decap_4 FILLER_8_668 ();
 sg13g2_fill_2 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_4 FILLER_8_721 ();
 sg13g2_fill_2 FILLER_8_725 ();
 sg13g2_fill_2 FILLER_8_732 ();
 sg13g2_fill_1 FILLER_8_734 ();
 sg13g2_decap_4 FILLER_8_743 ();
 sg13g2_decap_4 FILLER_8_764 ();
 sg13g2_fill_2 FILLER_8_768 ();
 sg13g2_fill_2 FILLER_8_778 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_fill_2 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_806 ();
 sg13g2_fill_2 FILLER_8_813 ();
 sg13g2_fill_1 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_fill_2 FILLER_8_850 ();
 sg13g2_fill_1 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_870 ();
 sg13g2_decap_8 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_8_884 ();
 sg13g2_decap_8 FILLER_8_891 ();
 sg13g2_decap_8 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_905 ();
 sg13g2_decap_8 FILLER_8_912 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_decap_8 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_933 ();
 sg13g2_decap_8 FILLER_8_940 ();
 sg13g2_decap_8 FILLER_8_947 ();
 sg13g2_decap_8 FILLER_8_954 ();
 sg13g2_decap_8 FILLER_8_961 ();
 sg13g2_decap_8 FILLER_8_968 ();
 sg13g2_decap_8 FILLER_8_975 ();
 sg13g2_decap_8 FILLER_8_982 ();
 sg13g2_decap_8 FILLER_8_989 ();
 sg13g2_decap_8 FILLER_8_996 ();
 sg13g2_decap_8 FILLER_8_1003 ();
 sg13g2_decap_8 FILLER_8_1010 ();
 sg13g2_decap_8 FILLER_8_1017 ();
 sg13g2_decap_4 FILLER_8_1024 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_2 FILLER_9_45 ();
 sg13g2_fill_1 FILLER_9_47 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_113 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_4 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_fill_2 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_fill_2 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_2 FILLER_9_435 ();
 sg13g2_decap_4 FILLER_9_441 ();
 sg13g2_fill_2 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_484 ();
 sg13g2_decap_4 FILLER_9_491 ();
 sg13g2_fill_1 FILLER_9_495 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_fill_2 FILLER_9_511 ();
 sg13g2_fill_1 FILLER_9_513 ();
 sg13g2_fill_1 FILLER_9_546 ();
 sg13g2_fill_1 FILLER_9_553 ();
 sg13g2_decap_4 FILLER_9_581 ();
 sg13g2_fill_2 FILLER_9_585 ();
 sg13g2_decap_4 FILLER_9_591 ();
 sg13g2_fill_2 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_601 ();
 sg13g2_fill_2 FILLER_9_608 ();
 sg13g2_fill_1 FILLER_9_610 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_fill_2 FILLER_9_651 ();
 sg13g2_fill_1 FILLER_9_658 ();
 sg13g2_decap_4 FILLER_9_666 ();
 sg13g2_fill_2 FILLER_9_670 ();
 sg13g2_fill_1 FILLER_9_684 ();
 sg13g2_fill_1 FILLER_9_699 ();
 sg13g2_fill_2 FILLER_9_708 ();
 sg13g2_decap_4 FILLER_9_715 ();
 sg13g2_fill_2 FILLER_9_719 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_fill_1 FILLER_9_746 ();
 sg13g2_fill_2 FILLER_9_767 ();
 sg13g2_fill_1 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_fill_2 FILLER_9_801 ();
 sg13g2_fill_1 FILLER_9_803 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_fill_2 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_832 ();
 sg13g2_decap_8 FILLER_9_839 ();
 sg13g2_fill_2 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_10_8 ();
 sg13g2_fill_1 FILLER_10_15 ();
 sg13g2_decap_8 FILLER_10_20 ();
 sg13g2_decap_8 FILLER_10_27 ();
 sg13g2_decap_4 FILLER_10_34 ();
 sg13g2_fill_1 FILLER_10_38 ();
 sg13g2_fill_1 FILLER_10_44 ();
 sg13g2_decap_4 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_58 ();
 sg13g2_decap_8 FILLER_10_69 ();
 sg13g2_fill_2 FILLER_10_76 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_decap_4 FILLER_10_83 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_decap_4 FILLER_10_155 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_172 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_decap_4 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_4 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_fill_1 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_fill_2 FILLER_10_373 ();
 sg13g2_decap_4 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_fill_1 FILLER_10_425 ();
 sg13g2_decap_8 FILLER_10_453 ();
 sg13g2_fill_2 FILLER_10_460 ();
 sg13g2_fill_2 FILLER_10_466 ();
 sg13g2_fill_2 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_482 ();
 sg13g2_fill_1 FILLER_10_489 ();
 sg13g2_decap_4 FILLER_10_508 ();
 sg13g2_fill_1 FILLER_10_512 ();
 sg13g2_fill_2 FILLER_10_531 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_fill_1 FILLER_10_581 ();
 sg13g2_fill_2 FILLER_10_610 ();
 sg13g2_fill_2 FILLER_10_617 ();
 sg13g2_decap_8 FILLER_10_635 ();
 sg13g2_decap_4 FILLER_10_642 ();
 sg13g2_fill_1 FILLER_10_646 ();
 sg13g2_decap_4 FILLER_10_675 ();
 sg13g2_fill_1 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_fill_1 FILLER_10_704 ();
 sg13g2_fill_2 FILLER_10_720 ();
 sg13g2_fill_1 FILLER_10_722 ();
 sg13g2_decap_4 FILLER_10_731 ();
 sg13g2_fill_2 FILLER_10_735 ();
 sg13g2_fill_2 FILLER_10_761 ();
 sg13g2_fill_2 FILLER_10_767 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_fill_2 FILLER_10_816 ();
 sg13g2_fill_1 FILLER_10_834 ();
 sg13g2_fill_2 FILLER_10_843 ();
 sg13g2_fill_1 FILLER_10_845 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_909 ();
 sg13g2_decap_8 FILLER_10_916 ();
 sg13g2_decap_8 FILLER_10_923 ();
 sg13g2_decap_8 FILLER_10_930 ();
 sg13g2_decap_8 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_951 ();
 sg13g2_decap_8 FILLER_10_958 ();
 sg13g2_decap_8 FILLER_10_965 ();
 sg13g2_decap_8 FILLER_10_972 ();
 sg13g2_decap_8 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_986 ();
 sg13g2_decap_8 FILLER_10_993 ();
 sg13g2_decap_8 FILLER_10_1000 ();
 sg13g2_decap_8 FILLER_10_1007 ();
 sg13g2_decap_8 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_fill_2 FILLER_11_67 ();
 sg13g2_decap_4 FILLER_11_79 ();
 sg13g2_fill_1 FILLER_11_83 ();
 sg13g2_decap_8 FILLER_11_90 ();
 sg13g2_decap_4 FILLER_11_115 ();
 sg13g2_decap_4 FILLER_11_133 ();
 sg13g2_decap_4 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_decap_4 FILLER_11_170 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_decap_4 FILLER_11_195 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_4 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_409 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_fill_2 FILLER_11_442 ();
 sg13g2_fill_2 FILLER_11_454 ();
 sg13g2_decap_8 FILLER_11_460 ();
 sg13g2_decap_4 FILLER_11_467 ();
 sg13g2_fill_1 FILLER_11_471 ();
 sg13g2_decap_8 FILLER_11_509 ();
 sg13g2_decap_4 FILLER_11_516 ();
 sg13g2_decap_4 FILLER_11_524 ();
 sg13g2_fill_1 FILLER_11_528 ();
 sg13g2_decap_4 FILLER_11_534 ();
 sg13g2_decap_4 FILLER_11_543 ();
 sg13g2_fill_2 FILLER_11_547 ();
 sg13g2_decap_8 FILLER_11_554 ();
 sg13g2_decap_8 FILLER_11_561 ();
 sg13g2_decap_8 FILLER_11_568 ();
 sg13g2_decap_4 FILLER_11_575 ();
 sg13g2_fill_1 FILLER_11_579 ();
 sg13g2_decap_8 FILLER_11_612 ();
 sg13g2_decap_8 FILLER_11_656 ();
 sg13g2_fill_2 FILLER_11_663 ();
 sg13g2_fill_1 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_671 ();
 sg13g2_decap_8 FILLER_11_678 ();
 sg13g2_decap_8 FILLER_11_685 ();
 sg13g2_fill_2 FILLER_11_692 ();
 sg13g2_fill_1 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_699 ();
 sg13g2_fill_1 FILLER_11_706 ();
 sg13g2_fill_2 FILLER_11_719 ();
 sg13g2_fill_1 FILLER_11_721 ();
 sg13g2_decap_4 FILLER_11_734 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_fill_2 FILLER_11_773 ();
 sg13g2_fill_1 FILLER_11_775 ();
 sg13g2_decap_8 FILLER_11_789 ();
 sg13g2_decap_4 FILLER_11_796 ();
 sg13g2_fill_1 FILLER_11_800 ();
 sg13g2_fill_2 FILLER_11_813 ();
 sg13g2_fill_1 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_834 ();
 sg13g2_decap_8 FILLER_11_841 ();
 sg13g2_decap_4 FILLER_11_848 ();
 sg13g2_fill_2 FILLER_11_862 ();
 sg13g2_fill_1 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_4 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_115 ();
 sg13g2_decap_4 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_4 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_201 ();
 sg13g2_decap_8 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_fill_1 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_4 FILLER_12_289 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_decap_4 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_332 ();
 sg13g2_decap_4 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_decap_8 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_12_436 ();
 sg13g2_decap_8 FILLER_12_442 ();
 sg13g2_fill_2 FILLER_12_449 ();
 sg13g2_decap_8 FILLER_12_478 ();
 sg13g2_fill_2 FILLER_12_485 ();
 sg13g2_fill_2 FILLER_12_491 ();
 sg13g2_fill_1 FILLER_12_493 ();
 sg13g2_decap_8 FILLER_12_498 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_fill_1 FILLER_12_568 ();
 sg13g2_decap_4 FILLER_12_579 ();
 sg13g2_fill_2 FILLER_12_583 ();
 sg13g2_decap_8 FILLER_12_589 ();
 sg13g2_fill_2 FILLER_12_596 ();
 sg13g2_fill_2 FILLER_12_610 ();
 sg13g2_fill_2 FILLER_12_620 ();
 sg13g2_fill_1 FILLER_12_622 ();
 sg13g2_fill_2 FILLER_12_627 ();
 sg13g2_fill_1 FILLER_12_633 ();
 sg13g2_decap_8 FILLER_12_638 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_4 FILLER_12_656 ();
 sg13g2_fill_1 FILLER_12_704 ();
 sg13g2_fill_1 FILLER_12_712 ();
 sg13g2_fill_1 FILLER_12_719 ();
 sg13g2_decap_8 FILLER_12_724 ();
 sg13g2_decap_4 FILLER_12_731 ();
 sg13g2_fill_1 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_762 ();
 sg13g2_fill_2 FILLER_12_769 ();
 sg13g2_fill_2 FILLER_12_794 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_fill_2 FILLER_12_816 ();
 sg13g2_decap_4 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_2 FILLER_12_861 ();
 sg13g2_fill_2 FILLER_12_876 ();
 sg13g2_decap_8 FILLER_12_891 ();
 sg13g2_decap_8 FILLER_12_898 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_decap_8 FILLER_12_912 ();
 sg13g2_decap_8 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_926 ();
 sg13g2_decap_8 FILLER_12_933 ();
 sg13g2_decap_8 FILLER_12_940 ();
 sg13g2_decap_8 FILLER_12_947 ();
 sg13g2_decap_8 FILLER_12_954 ();
 sg13g2_decap_8 FILLER_12_961 ();
 sg13g2_decap_8 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_975 ();
 sg13g2_decap_8 FILLER_12_982 ();
 sg13g2_decap_8 FILLER_12_989 ();
 sg13g2_decap_8 FILLER_12_996 ();
 sg13g2_decap_8 FILLER_12_1003 ();
 sg13g2_decap_8 FILLER_12_1010 ();
 sg13g2_decap_8 FILLER_12_1017 ();
 sg13g2_decap_4 FILLER_12_1024 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_4 FILLER_13_4 ();
 sg13g2_fill_2 FILLER_13_8 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_decap_8 FILLER_13_44 ();
 sg13g2_decap_4 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_55 ();
 sg13g2_decap_8 FILLER_13_61 ();
 sg13g2_decap_8 FILLER_13_68 ();
 sg13g2_decap_8 FILLER_13_75 ();
 sg13g2_fill_1 FILLER_13_82 ();
 sg13g2_fill_1 FILLER_13_114 ();
 sg13g2_decap_4 FILLER_13_125 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_4 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_170 ();
 sg13g2_decap_4 FILLER_13_177 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_decap_4 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_decap_4 FILLER_13_328 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_2 FILLER_13_355 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_4 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_13_406 ();
 sg13g2_fill_2 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_453 ();
 sg13g2_decap_8 FILLER_13_460 ();
 sg13g2_decap_8 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_fill_2 FILLER_13_492 ();
 sg13g2_fill_1 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_505 ();
 sg13g2_decap_8 FILLER_13_512 ();
 sg13g2_decap_8 FILLER_13_519 ();
 sg13g2_decap_4 FILLER_13_526 ();
 sg13g2_fill_2 FILLER_13_530 ();
 sg13g2_fill_2 FILLER_13_542 ();
 sg13g2_fill_1 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_4 FILLER_13_586 ();
 sg13g2_fill_2 FILLER_13_590 ();
 sg13g2_decap_8 FILLER_13_617 ();
 sg13g2_fill_2 FILLER_13_624 ();
 sg13g2_fill_1 FILLER_13_626 ();
 sg13g2_fill_2 FILLER_13_637 ();
 sg13g2_fill_1 FILLER_13_639 ();
 sg13g2_fill_1 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_4 FILLER_13_684 ();
 sg13g2_fill_2 FILLER_13_688 ();
 sg13g2_fill_2 FILLER_13_698 ();
 sg13g2_decap_4 FILLER_13_704 ();
 sg13g2_fill_1 FILLER_13_708 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_fill_2 FILLER_13_728 ();
 sg13g2_fill_2 FILLER_13_740 ();
 sg13g2_fill_2 FILLER_13_755 ();
 sg13g2_decap_8 FILLER_13_766 ();
 sg13g2_fill_2 FILLER_13_773 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_fill_1 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_fill_2 FILLER_13_837 ();
 sg13g2_fill_1 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_848 ();
 sg13g2_decap_8 FILLER_13_855 ();
 sg13g2_decap_8 FILLER_13_862 ();
 sg13g2_fill_2 FILLER_13_869 ();
 sg13g2_fill_2 FILLER_13_883 ();
 sg13g2_fill_1 FILLER_13_885 ();
 sg13g2_decap_8 FILLER_13_891 ();
 sg13g2_decap_8 FILLER_13_898 ();
 sg13g2_decap_8 FILLER_13_905 ();
 sg13g2_decap_8 FILLER_13_912 ();
 sg13g2_decap_8 FILLER_13_919 ();
 sg13g2_decap_8 FILLER_13_926 ();
 sg13g2_decap_8 FILLER_13_933 ();
 sg13g2_decap_8 FILLER_13_940 ();
 sg13g2_decap_8 FILLER_13_947 ();
 sg13g2_decap_8 FILLER_13_954 ();
 sg13g2_decap_8 FILLER_13_961 ();
 sg13g2_decap_8 FILLER_13_968 ();
 sg13g2_decap_8 FILLER_13_975 ();
 sg13g2_decap_8 FILLER_13_982 ();
 sg13g2_decap_8 FILLER_13_989 ();
 sg13g2_decap_8 FILLER_13_996 ();
 sg13g2_decap_8 FILLER_13_1003 ();
 sg13g2_decap_8 FILLER_13_1010 ();
 sg13g2_decap_8 FILLER_13_1017 ();
 sg13g2_decap_4 FILLER_13_1024 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_4 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_8 ();
 sg13g2_fill_2 FILLER_14_17 ();
 sg13g2_fill_1 FILLER_14_19 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_decap_8 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_86 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_decap_4 FILLER_14_96 ();
 sg13g2_decap_8 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_111 ();
 sg13g2_decap_4 FILLER_14_119 ();
 sg13g2_decap_4 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_decap_4 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_decap_4 FILLER_14_409 ();
 sg13g2_fill_2 FILLER_14_413 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_14_439 ();
 sg13g2_fill_2 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_fill_2 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_4 FILLER_14_591 ();
 sg13g2_fill_1 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_615 ();
 sg13g2_decap_8 FILLER_14_622 ();
 sg13g2_fill_2 FILLER_14_629 ();
 sg13g2_fill_1 FILLER_14_645 ();
 sg13g2_fill_2 FILLER_14_674 ();
 sg13g2_fill_1 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_706 ();
 sg13g2_decap_8 FILLER_14_713 ();
 sg13g2_fill_2 FILLER_14_720 ();
 sg13g2_fill_1 FILLER_14_722 ();
 sg13g2_decap_4 FILLER_14_757 ();
 sg13g2_fill_2 FILLER_14_761 ();
 sg13g2_fill_2 FILLER_14_769 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_4 FILLER_14_798 ();
 sg13g2_fill_2 FILLER_14_810 ();
 sg13g2_fill_1 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_825 ();
 sg13g2_fill_2 FILLER_14_832 ();
 sg13g2_fill_1 FILLER_14_834 ();
 sg13g2_fill_2 FILLER_14_862 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_8 FILLER_14_910 ();
 sg13g2_decap_8 FILLER_14_917 ();
 sg13g2_decap_8 FILLER_14_924 ();
 sg13g2_decap_8 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_decap_8 FILLER_14_945 ();
 sg13g2_decap_8 FILLER_14_952 ();
 sg13g2_decap_8 FILLER_14_959 ();
 sg13g2_decap_8 FILLER_14_966 ();
 sg13g2_decap_8 FILLER_14_973 ();
 sg13g2_decap_8 FILLER_14_980 ();
 sg13g2_decap_8 FILLER_14_987 ();
 sg13g2_decap_8 FILLER_14_994 ();
 sg13g2_decap_8 FILLER_14_1001 ();
 sg13g2_decap_8 FILLER_14_1008 ();
 sg13g2_decap_8 FILLER_14_1015 ();
 sg13g2_decap_8 FILLER_14_1022 ();
 sg13g2_decap_4 FILLER_15_4 ();
 sg13g2_decap_4 FILLER_15_45 ();
 sg13g2_fill_2 FILLER_15_116 ();
 sg13g2_fill_1 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_4 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_4 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_354 ();
 sg13g2_decap_4 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_4 FILLER_15_406 ();
 sg13g2_fill_2 FILLER_15_410 ();
 sg13g2_fill_2 FILLER_15_426 ();
 sg13g2_fill_1 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_fill_1 FILLER_15_473 ();
 sg13g2_decap_4 FILLER_15_478 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_fill_1 FILLER_15_506 ();
 sg13g2_fill_2 FILLER_15_511 ();
 sg13g2_fill_1 FILLER_15_513 ();
 sg13g2_decap_4 FILLER_15_518 ();
 sg13g2_fill_2 FILLER_15_522 ();
 sg13g2_decap_4 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_4 FILLER_15_550 ();
 sg13g2_decap_4 FILLER_15_558 ();
 sg13g2_decap_8 FILLER_15_580 ();
 sg13g2_fill_1 FILLER_15_587 ();
 sg13g2_fill_1 FILLER_15_599 ();
 sg13g2_fill_2 FILLER_15_615 ();
 sg13g2_fill_1 FILLER_15_617 ();
 sg13g2_decap_4 FILLER_15_646 ();
 sg13g2_fill_1 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_fill_1 FILLER_15_690 ();
 sg13g2_decap_4 FILLER_15_696 ();
 sg13g2_decap_4 FILLER_15_708 ();
 sg13g2_decap_4 FILLER_15_748 ();
 sg13g2_fill_2 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_758 ();
 sg13g2_decap_8 FILLER_15_765 ();
 sg13g2_decap_4 FILLER_15_772 ();
 sg13g2_fill_1 FILLER_15_776 ();
 sg13g2_decap_4 FILLER_15_785 ();
 sg13g2_fill_2 FILLER_15_789 ();
 sg13g2_decap_8 FILLER_15_797 ();
 sg13g2_fill_1 FILLER_15_804 ();
 sg13g2_fill_2 FILLER_15_818 ();
 sg13g2_decap_8 FILLER_15_828 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_fill_2 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_4 FILLER_15_868 ();
 sg13g2_fill_2 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_891 ();
 sg13g2_decap_8 FILLER_15_898 ();
 sg13g2_decap_8 FILLER_15_905 ();
 sg13g2_decap_8 FILLER_15_912 ();
 sg13g2_decap_8 FILLER_15_919 ();
 sg13g2_decap_8 FILLER_15_926 ();
 sg13g2_decap_8 FILLER_15_933 ();
 sg13g2_decap_8 FILLER_15_940 ();
 sg13g2_decap_8 FILLER_15_947 ();
 sg13g2_decap_8 FILLER_15_954 ();
 sg13g2_decap_8 FILLER_15_961 ();
 sg13g2_decap_8 FILLER_15_968 ();
 sg13g2_decap_8 FILLER_15_975 ();
 sg13g2_decap_8 FILLER_15_982 ();
 sg13g2_decap_8 FILLER_15_989 ();
 sg13g2_decap_8 FILLER_15_996 ();
 sg13g2_decap_8 FILLER_15_1003 ();
 sg13g2_decap_8 FILLER_15_1010 ();
 sg13g2_decap_8 FILLER_15_1017 ();
 sg13g2_decap_4 FILLER_15_1024 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_4 FILLER_16_4 ();
 sg13g2_decap_4 FILLER_16_45 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_85 ();
 sg13g2_decap_8 FILLER_16_97 ();
 sg13g2_decap_4 FILLER_16_104 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_148 ();
 sg13g2_decap_8 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_fill_2 FILLER_16_387 ();
 sg13g2_fill_1 FILLER_16_389 ();
 sg13g2_fill_1 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_fill_2 FILLER_16_450 ();
 sg13g2_fill_1 FILLER_16_452 ();
 sg13g2_fill_2 FILLER_16_480 ();
 sg13g2_fill_1 FILLER_16_482 ();
 sg13g2_decap_4 FILLER_16_487 ();
 sg13g2_fill_2 FILLER_16_516 ();
 sg13g2_fill_1 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_4 FILLER_16_589 ();
 sg13g2_fill_2 FILLER_16_593 ();
 sg13g2_fill_2 FILLER_16_607 ();
 sg13g2_decap_4 FILLER_16_617 ();
 sg13g2_fill_2 FILLER_16_621 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_4 FILLER_16_653 ();
 sg13g2_fill_2 FILLER_16_657 ();
 sg13g2_fill_1 FILLER_16_664 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_fill_2 FILLER_16_679 ();
 sg13g2_fill_1 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_fill_1 FILLER_16_718 ();
 sg13g2_fill_2 FILLER_16_733 ();
 sg13g2_fill_1 FILLER_16_746 ();
 sg13g2_decap_4 FILLER_16_762 ();
 sg13g2_decap_8 FILLER_16_778 ();
 sg13g2_fill_2 FILLER_16_785 ();
 sg13g2_fill_1 FILLER_16_787 ();
 sg13g2_decap_4 FILLER_16_804 ();
 sg13g2_fill_1 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_fill_1 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_fill_2 FILLER_16_868 ();
 sg13g2_fill_1 FILLER_16_870 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_decap_8 FILLER_17_4 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_decap_4 FILLER_17_17 ();
 sg13g2_decap_8 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_120 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_decap_4 FILLER_17_144 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_174 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_376 ();
 sg13g2_fill_1 FILLER_17_378 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_1 FILLER_17_400 ();
 sg13g2_decap_4 FILLER_17_432 ();
 sg13g2_decap_8 FILLER_17_440 ();
 sg13g2_decap_8 FILLER_17_451 ();
 sg13g2_decap_4 FILLER_17_458 ();
 sg13g2_fill_1 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_fill_2 FILLER_17_549 ();
 sg13g2_fill_2 FILLER_17_564 ();
 sg13g2_fill_2 FILLER_17_571 ();
 sg13g2_fill_1 FILLER_17_573 ();
 sg13g2_decap_8 FILLER_17_579 ();
 sg13g2_decap_4 FILLER_17_586 ();
 sg13g2_fill_1 FILLER_17_590 ();
 sg13g2_decap_8 FILLER_17_619 ();
 sg13g2_decap_8 FILLER_17_626 ();
 sg13g2_fill_2 FILLER_17_633 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_737 ();
 sg13g2_decap_8 FILLER_17_744 ();
 sg13g2_decap_8 FILLER_17_751 ();
 sg13g2_fill_2 FILLER_17_758 ();
 sg13g2_fill_1 FILLER_17_760 ();
 sg13g2_fill_2 FILLER_17_766 ();
 sg13g2_fill_1 FILLER_17_768 ();
 sg13g2_decap_4 FILLER_17_779 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_4 FILLER_17_836 ();
 sg13g2_fill_1 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_860 ();
 sg13g2_decap_4 FILLER_17_867 ();
 sg13g2_fill_1 FILLER_17_871 ();
 sg13g2_decap_8 FILLER_17_898 ();
 sg13g2_decap_8 FILLER_17_905 ();
 sg13g2_decap_8 FILLER_17_912 ();
 sg13g2_decap_8 FILLER_17_919 ();
 sg13g2_decap_8 FILLER_17_926 ();
 sg13g2_decap_8 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_940 ();
 sg13g2_decap_8 FILLER_17_947 ();
 sg13g2_decap_8 FILLER_17_954 ();
 sg13g2_decap_8 FILLER_17_961 ();
 sg13g2_decap_8 FILLER_17_968 ();
 sg13g2_decap_8 FILLER_17_975 ();
 sg13g2_decap_8 FILLER_17_982 ();
 sg13g2_decap_8 FILLER_17_989 ();
 sg13g2_decap_8 FILLER_17_996 ();
 sg13g2_decap_8 FILLER_17_1003 ();
 sg13g2_decap_8 FILLER_17_1010 ();
 sg13g2_decap_8 FILLER_17_1017 ();
 sg13g2_decap_4 FILLER_17_1024 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_decap_8 FILLER_18_37 ();
 sg13g2_fill_2 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_4 FILLER_18_195 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_4 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_decap_4 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_fill_1 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_458 ();
 sg13g2_fill_1 FILLER_18_460 ();
 sg13g2_fill_2 FILLER_18_465 ();
 sg13g2_fill_1 FILLER_18_467 ();
 sg13g2_fill_2 FILLER_18_472 ();
 sg13g2_decap_8 FILLER_18_478 ();
 sg13g2_decap_4 FILLER_18_491 ();
 sg13g2_fill_1 FILLER_18_495 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_4 FILLER_18_508 ();
 sg13g2_fill_1 FILLER_18_512 ();
 sg13g2_decap_8 FILLER_18_521 ();
 sg13g2_fill_2 FILLER_18_528 ();
 sg13g2_fill_1 FILLER_18_534 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_fill_2 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_583 ();
 sg13g2_decap_4 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_614 ();
 sg13g2_decap_4 FILLER_18_647 ();
 sg13g2_fill_2 FILLER_18_651 ();
 sg13g2_fill_2 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_669 ();
 sg13g2_fill_1 FILLER_18_688 ();
 sg13g2_fill_2 FILLER_18_694 ();
 sg13g2_fill_1 FILLER_18_696 ();
 sg13g2_decap_8 FILLER_18_705 ();
 sg13g2_decap_8 FILLER_18_712 ();
 sg13g2_fill_2 FILLER_18_719 ();
 sg13g2_decap_8 FILLER_18_741 ();
 sg13g2_fill_1 FILLER_18_748 ();
 sg13g2_decap_4 FILLER_18_755 ();
 sg13g2_fill_1 FILLER_18_759 ();
 sg13g2_fill_2 FILLER_18_765 ();
 sg13g2_decap_4 FILLER_18_780 ();
 sg13g2_fill_1 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_4 FILLER_18_799 ();
 sg13g2_fill_2 FILLER_18_803 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_fill_2 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_863 ();
 sg13g2_decap_4 FILLER_18_870 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_decap_8 FILLER_18_912 ();
 sg13g2_decap_8 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_decap_8 FILLER_18_954 ();
 sg13g2_decap_8 FILLER_18_961 ();
 sg13g2_decap_8 FILLER_18_968 ();
 sg13g2_decap_8 FILLER_18_975 ();
 sg13g2_decap_8 FILLER_18_982 ();
 sg13g2_decap_8 FILLER_18_989 ();
 sg13g2_decap_8 FILLER_18_996 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1010 ();
 sg13g2_decap_8 FILLER_18_1017 ();
 sg13g2_decap_4 FILLER_18_1024 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_9 ();
 sg13g2_fill_1 FILLER_19_16 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_4 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_72 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_decap_4 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_decap_4 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_282 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_decap_4 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_decap_4 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_2 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_19_410 ();
 sg13g2_decap_4 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_425 ();
 sg13g2_decap_4 FILLER_19_445 ();
 sg13g2_fill_2 FILLER_19_476 ();
 sg13g2_fill_1 FILLER_19_478 ();
 sg13g2_decap_8 FILLER_19_493 ();
 sg13g2_decap_8 FILLER_19_500 ();
 sg13g2_decap_4 FILLER_19_507 ();
 sg13g2_fill_1 FILLER_19_511 ();
 sg13g2_fill_2 FILLER_19_522 ();
 sg13g2_fill_1 FILLER_19_524 ();
 sg13g2_decap_8 FILLER_19_552 ();
 sg13g2_fill_2 FILLER_19_559 ();
 sg13g2_decap_4 FILLER_19_565 ();
 sg13g2_fill_2 FILLER_19_569 ();
 sg13g2_decap_8 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_587 ();
 sg13g2_decap_8 FILLER_19_612 ();
 sg13g2_fill_1 FILLER_19_619 ();
 sg13g2_decap_8 FILLER_19_624 ();
 sg13g2_decap_8 FILLER_19_631 ();
 sg13g2_decap_8 FILLER_19_638 ();
 sg13g2_fill_2 FILLER_19_645 ();
 sg13g2_fill_1 FILLER_19_647 ();
 sg13g2_fill_2 FILLER_19_653 ();
 sg13g2_fill_1 FILLER_19_655 ();
 sg13g2_decap_4 FILLER_19_665 ();
 sg13g2_fill_2 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_4 FILLER_19_711 ();
 sg13g2_fill_1 FILLER_19_715 ();
 sg13g2_decap_8 FILLER_19_744 ();
 sg13g2_fill_2 FILLER_19_759 ();
 sg13g2_fill_1 FILLER_19_761 ();
 sg13g2_decap_4 FILLER_19_772 ();
 sg13g2_fill_2 FILLER_19_776 ();
 sg13g2_decap_8 FILLER_19_792 ();
 sg13g2_fill_2 FILLER_19_819 ();
 sg13g2_fill_1 FILLER_19_821 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_fill_1 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_855 ();
 sg13g2_decap_8 FILLER_19_862 ();
 sg13g2_decap_8 FILLER_19_869 ();
 sg13g2_decap_4 FILLER_19_876 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_8 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_930 ();
 sg13g2_decap_8 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_944 ();
 sg13g2_decap_8 FILLER_19_951 ();
 sg13g2_decap_8 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_decap_8 FILLER_19_1000 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_4 FILLER_19_1021 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_fill_1 FILLER_20_20 ();
 sg13g2_fill_1 FILLER_20_58 ();
 sg13g2_decap_4 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_decap_4 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_fill_1 FILLER_20_418 ();
 sg13g2_fill_1 FILLER_20_424 ();
 sg13g2_decap_4 FILLER_20_435 ();
 sg13g2_fill_2 FILLER_20_439 ();
 sg13g2_fill_2 FILLER_20_451 ();
 sg13g2_fill_1 FILLER_20_453 ();
 sg13g2_decap_8 FILLER_20_458 ();
 sg13g2_decap_8 FILLER_20_465 ();
 sg13g2_decap_4 FILLER_20_472 ();
 sg13g2_fill_1 FILLER_20_476 ();
 sg13g2_fill_1 FILLER_20_508 ();
 sg13g2_decap_8 FILLER_20_519 ();
 sg13g2_fill_1 FILLER_20_526 ();
 sg13g2_fill_2 FILLER_20_531 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_decap_4 FILLER_20_565 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_decap_8 FILLER_20_598 ();
 sg13g2_decap_4 FILLER_20_605 ();
 sg13g2_fill_2 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_4 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_fill_2 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_4 FILLER_20_713 ();
 sg13g2_fill_1 FILLER_20_727 ();
 sg13g2_decap_4 FILLER_20_735 ();
 sg13g2_fill_2 FILLER_20_739 ();
 sg13g2_decap_8 FILLER_20_745 ();
 sg13g2_fill_1 FILLER_20_752 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_787 ();
 sg13g2_decap_8 FILLER_20_794 ();
 sg13g2_decap_4 FILLER_20_801 ();
 sg13g2_decap_4 FILLER_20_815 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_852 ();
 sg13g2_fill_2 FILLER_20_859 ();
 sg13g2_decap_8 FILLER_20_906 ();
 sg13g2_decap_8 FILLER_20_913 ();
 sg13g2_decap_8 FILLER_20_920 ();
 sg13g2_decap_8 FILLER_20_927 ();
 sg13g2_decap_8 FILLER_20_934 ();
 sg13g2_decap_8 FILLER_20_941 ();
 sg13g2_decap_8 FILLER_20_948 ();
 sg13g2_decap_8 FILLER_20_955 ();
 sg13g2_decap_8 FILLER_20_962 ();
 sg13g2_decap_8 FILLER_20_969 ();
 sg13g2_decap_8 FILLER_20_976 ();
 sg13g2_decap_8 FILLER_20_983 ();
 sg13g2_decap_8 FILLER_20_990 ();
 sg13g2_decap_8 FILLER_20_997 ();
 sg13g2_decap_8 FILLER_20_1004 ();
 sg13g2_decap_8 FILLER_20_1011 ();
 sg13g2_decap_8 FILLER_20_1018 ();
 sg13g2_decap_4 FILLER_20_1025 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_30 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_decap_8 FILLER_21_76 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_4 FILLER_21_170 ();
 sg13g2_decap_4 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_4 FILLER_21_276 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_21_457 ();
 sg13g2_fill_1 FILLER_21_464 ();
 sg13g2_fill_1 FILLER_21_489 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_fill_1 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_decap_8 FILLER_21_556 ();
 sg13g2_decap_4 FILLER_21_563 ();
 sg13g2_fill_1 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_592 ();
 sg13g2_fill_1 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_fill_2 FILLER_21_645 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_fill_2 FILLER_21_679 ();
 sg13g2_decap_4 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_701 ();
 sg13g2_decap_8 FILLER_21_737 ();
 sg13g2_decap_4 FILLER_21_744 ();
 sg13g2_fill_1 FILLER_21_748 ();
 sg13g2_fill_2 FILLER_21_774 ();
 sg13g2_fill_1 FILLER_21_776 ();
 sg13g2_decap_4 FILLER_21_793 ();
 sg13g2_fill_1 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_4 FILLER_21_830 ();
 sg13g2_fill_1 FILLER_21_834 ();
 sg13g2_decap_8 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_21_865 ();
 sg13g2_fill_2 FILLER_21_872 ();
 sg13g2_fill_1 FILLER_21_874 ();
 sg13g2_decap_8 FILLER_21_901 ();
 sg13g2_decap_8 FILLER_21_908 ();
 sg13g2_decap_8 FILLER_21_915 ();
 sg13g2_decap_8 FILLER_21_922 ();
 sg13g2_decap_8 FILLER_21_929 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_950 ();
 sg13g2_decap_8 FILLER_21_957 ();
 sg13g2_decap_8 FILLER_21_964 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_decap_8 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_985 ();
 sg13g2_decap_8 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_999 ();
 sg13g2_decap_8 FILLER_21_1006 ();
 sg13g2_decap_8 FILLER_21_1013 ();
 sg13g2_decap_8 FILLER_21_1020 ();
 sg13g2_fill_2 FILLER_21_1027 ();
 sg13g2_decap_4 FILLER_22_8 ();
 sg13g2_fill_1 FILLER_22_12 ();
 sg13g2_fill_2 FILLER_22_17 ();
 sg13g2_fill_1 FILLER_22_19 ();
 sg13g2_decap_8 FILLER_22_47 ();
 sg13g2_decap_4 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_4 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_4 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_308 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_339 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_decap_4 FILLER_22_393 ();
 sg13g2_fill_1 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_402 ();
 sg13g2_decap_4 FILLER_22_410 ();
 sg13g2_fill_1 FILLER_22_414 ();
 sg13g2_fill_2 FILLER_22_420 ();
 sg13g2_fill_1 FILLER_22_422 ();
 sg13g2_fill_2 FILLER_22_448 ();
 sg13g2_fill_1 FILLER_22_450 ();
 sg13g2_fill_1 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_505 ();
 sg13g2_decap_8 FILLER_22_512 ();
 sg13g2_decap_4 FILLER_22_519 ();
 sg13g2_decap_4 FILLER_22_527 ();
 sg13g2_decap_8 FILLER_22_562 ();
 sg13g2_decap_4 FILLER_22_569 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_600 ();
 sg13g2_fill_1 FILLER_22_607 ();
 sg13g2_fill_1 FILLER_22_621 ();
 sg13g2_decap_8 FILLER_22_695 ();
 sg13g2_decap_4 FILLER_22_702 ();
 sg13g2_fill_2 FILLER_22_706 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_4 FILLER_22_747 ();
 sg13g2_fill_1 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_fill_2 FILLER_22_797 ();
 sg13g2_decap_8 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_824 ();
 sg13g2_fill_2 FILLER_22_831 ();
 sg13g2_decap_8 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_22_862 ();
 sg13g2_fill_2 FILLER_22_869 ();
 sg13g2_decap_8 FILLER_22_897 ();
 sg13g2_decap_8 FILLER_22_904 ();
 sg13g2_decap_8 FILLER_22_911 ();
 sg13g2_decap_8 FILLER_22_918 ();
 sg13g2_decap_8 FILLER_22_925 ();
 sg13g2_decap_8 FILLER_22_932 ();
 sg13g2_decap_8 FILLER_22_939 ();
 sg13g2_decap_8 FILLER_22_946 ();
 sg13g2_decap_8 FILLER_22_953 ();
 sg13g2_decap_8 FILLER_22_960 ();
 sg13g2_decap_8 FILLER_22_967 ();
 sg13g2_decap_8 FILLER_22_974 ();
 sg13g2_decap_8 FILLER_22_981 ();
 sg13g2_decap_8 FILLER_22_988 ();
 sg13g2_decap_8 FILLER_22_995 ();
 sg13g2_decap_8 FILLER_22_1002 ();
 sg13g2_decap_8 FILLER_22_1009 ();
 sg13g2_decap_8 FILLER_22_1016 ();
 sg13g2_decap_4 FILLER_22_1023 ();
 sg13g2_fill_2 FILLER_22_1027 ();
 sg13g2_fill_1 FILLER_23_31 ();
 sg13g2_decap_4 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_fill_2 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_4 FILLER_23_192 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_decap_8 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_4 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_23_440 ();
 sg13g2_decap_8 FILLER_23_454 ();
 sg13g2_fill_2 FILLER_23_461 ();
 sg13g2_decap_4 FILLER_23_467 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_4 FILLER_23_487 ();
 sg13g2_fill_2 FILLER_23_491 ();
 sg13g2_fill_1 FILLER_23_510 ();
 sg13g2_fill_2 FILLER_23_538 ();
 sg13g2_decap_8 FILLER_23_544 ();
 sg13g2_fill_2 FILLER_23_551 ();
 sg13g2_fill_1 FILLER_23_553 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_4 FILLER_23_578 ();
 sg13g2_decap_4 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_8 FILLER_23_640 ();
 sg13g2_decap_8 FILLER_23_647 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_fill_1 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_fill_2 FILLER_23_690 ();
 sg13g2_fill_1 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_736 ();
 sg13g2_fill_2 FILLER_23_743 ();
 sg13g2_fill_1 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_771 ();
 sg13g2_fill_2 FILLER_23_778 ();
 sg13g2_fill_2 FILLER_23_796 ();
 sg13g2_fill_1 FILLER_23_798 ();
 sg13g2_fill_2 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_decap_8 FILLER_23_820 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_fill_1 FILLER_23_859 ();
 sg13g2_decap_8 FILLER_23_895 ();
 sg13g2_decap_8 FILLER_23_902 ();
 sg13g2_decap_8 FILLER_23_909 ();
 sg13g2_decap_8 FILLER_23_916 ();
 sg13g2_decap_8 FILLER_23_923 ();
 sg13g2_decap_8 FILLER_23_930 ();
 sg13g2_decap_8 FILLER_23_937 ();
 sg13g2_decap_8 FILLER_23_944 ();
 sg13g2_decap_8 FILLER_23_951 ();
 sg13g2_decap_8 FILLER_23_958 ();
 sg13g2_decap_8 FILLER_23_965 ();
 sg13g2_decap_8 FILLER_23_972 ();
 sg13g2_decap_8 FILLER_23_979 ();
 sg13g2_decap_8 FILLER_23_986 ();
 sg13g2_decap_8 FILLER_23_993 ();
 sg13g2_decap_8 FILLER_23_1000 ();
 sg13g2_decap_8 FILLER_23_1007 ();
 sg13g2_decap_8 FILLER_23_1014 ();
 sg13g2_decap_8 FILLER_23_1021 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_9 ();
 sg13g2_decap_8 FILLER_24_36 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_decap_8 FILLER_24_71 ();
 sg13g2_decap_4 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_4 FILLER_24_100 ();
 sg13g2_decap_4 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_decap_4 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_4 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_4 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_405 ();
 sg13g2_fill_2 FILLER_24_449 ();
 sg13g2_fill_1 FILLER_24_451 ();
 sg13g2_decap_4 FILLER_24_479 ();
 sg13g2_fill_2 FILLER_24_483 ();
 sg13g2_decap_4 FILLER_24_489 ();
 sg13g2_decap_4 FILLER_24_497 ();
 sg13g2_fill_2 FILLER_24_501 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_520 ();
 sg13g2_decap_4 FILLER_24_527 ();
 sg13g2_fill_1 FILLER_24_531 ();
 sg13g2_decap_8 FILLER_24_590 ();
 sg13g2_decap_8 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_612 ();
 sg13g2_decap_8 FILLER_24_619 ();
 sg13g2_decap_8 FILLER_24_626 ();
 sg13g2_decap_8 FILLER_24_633 ();
 sg13g2_decap_4 FILLER_24_640 ();
 sg13g2_fill_2 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_4 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_687 ();
 sg13g2_decap_8 FILLER_24_694 ();
 sg13g2_fill_2 FILLER_24_701 ();
 sg13g2_fill_1 FILLER_24_703 ();
 sg13g2_fill_2 FILLER_24_709 ();
 sg13g2_fill_1 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_fill_1 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_4 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_4 FILLER_24_831 ();
 sg13g2_fill_2 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_4 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_885 ();
 sg13g2_decap_8 FILLER_24_892 ();
 sg13g2_decap_8 FILLER_24_899 ();
 sg13g2_decap_8 FILLER_24_906 ();
 sg13g2_decap_8 FILLER_24_913 ();
 sg13g2_decap_8 FILLER_24_920 ();
 sg13g2_decap_8 FILLER_24_927 ();
 sg13g2_decap_8 FILLER_24_934 ();
 sg13g2_decap_8 FILLER_24_941 ();
 sg13g2_decap_8 FILLER_24_948 ();
 sg13g2_decap_8 FILLER_24_955 ();
 sg13g2_decap_8 FILLER_24_962 ();
 sg13g2_decap_8 FILLER_24_969 ();
 sg13g2_decap_8 FILLER_24_976 ();
 sg13g2_decap_8 FILLER_24_983 ();
 sg13g2_decap_8 FILLER_24_990 ();
 sg13g2_decap_8 FILLER_24_997 ();
 sg13g2_decap_8 FILLER_24_1004 ();
 sg13g2_decap_8 FILLER_24_1011 ();
 sg13g2_decap_8 FILLER_24_1018 ();
 sg13g2_decap_4 FILLER_24_1025 ();
 sg13g2_decap_4 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_73 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_4 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_decap_4 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_4 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_4 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_fill_2 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_436 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_decap_8 FILLER_25_450 ();
 sg13g2_decap_8 FILLER_25_461 ();
 sg13g2_decap_8 FILLER_25_468 ();
 sg13g2_fill_2 FILLER_25_475 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_fill_1 FILLER_25_516 ();
 sg13g2_fill_1 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_decap_8 FILLER_25_534 ();
 sg13g2_decap_8 FILLER_25_545 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_4 FILLER_25_566 ();
 sg13g2_fill_2 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_fill_1 FILLER_25_654 ();
 sg13g2_fill_1 FILLER_25_663 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_684 ();
 sg13g2_fill_1 FILLER_25_691 ();
 sg13g2_fill_2 FILLER_25_700 ();
 sg13g2_fill_1 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_4 FILLER_25_749 ();
 sg13g2_fill_1 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_759 ();
 sg13g2_decap_8 FILLER_25_766 ();
 sg13g2_decap_4 FILLER_25_773 ();
 sg13g2_fill_1 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_fill_1 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_25_865 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_decap_8 FILLER_25_893 ();
 sg13g2_decap_8 FILLER_25_900 ();
 sg13g2_decap_8 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_914 ();
 sg13g2_decap_8 FILLER_25_921 ();
 sg13g2_decap_8 FILLER_25_928 ();
 sg13g2_decap_8 FILLER_25_935 ();
 sg13g2_decap_8 FILLER_25_942 ();
 sg13g2_decap_8 FILLER_25_949 ();
 sg13g2_decap_8 FILLER_25_956 ();
 sg13g2_decap_8 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_970 ();
 sg13g2_decap_8 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_984 ();
 sg13g2_decap_8 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_998 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_8 FILLER_25_1012 ();
 sg13g2_decap_8 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_fill_1 FILLER_26_13 ();
 sg13g2_fill_2 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_24 ();
 sg13g2_decap_8 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_decap_4 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_232 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_4 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_4 FILLER_26_473 ();
 sg13g2_decap_4 FILLER_26_491 ();
 sg13g2_fill_2 FILLER_26_495 ();
 sg13g2_decap_4 FILLER_26_545 ();
 sg13g2_fill_1 FILLER_26_549 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_fill_1 FILLER_26_567 ();
 sg13g2_decap_4 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_610 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_fill_1 FILLER_26_668 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_fill_2 FILLER_26_686 ();
 sg13g2_fill_2 FILLER_26_697 ();
 sg13g2_fill_2 FILLER_26_703 ();
 sg13g2_decap_8 FILLER_26_710 ();
 sg13g2_decap_4 FILLER_26_717 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_4 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_4 FILLER_26_785 ();
 sg13g2_fill_2 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_decap_8 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_853 ();
 sg13g2_decap_8 FILLER_26_860 ();
 sg13g2_decap_8 FILLER_26_867 ();
 sg13g2_decap_8 FILLER_26_874 ();
 sg13g2_decap_8 FILLER_26_881 ();
 sg13g2_decap_8 FILLER_26_888 ();
 sg13g2_decap_8 FILLER_26_895 ();
 sg13g2_decap_8 FILLER_26_902 ();
 sg13g2_decap_8 FILLER_26_909 ();
 sg13g2_decap_8 FILLER_26_916 ();
 sg13g2_decap_8 FILLER_26_923 ();
 sg13g2_decap_8 FILLER_26_930 ();
 sg13g2_decap_8 FILLER_26_937 ();
 sg13g2_decap_8 FILLER_26_944 ();
 sg13g2_decap_8 FILLER_26_951 ();
 sg13g2_decap_8 FILLER_26_958 ();
 sg13g2_decap_8 FILLER_26_965 ();
 sg13g2_decap_8 FILLER_26_972 ();
 sg13g2_decap_8 FILLER_26_979 ();
 sg13g2_decap_8 FILLER_26_986 ();
 sg13g2_decap_8 FILLER_26_993 ();
 sg13g2_decap_8 FILLER_26_1000 ();
 sg13g2_decap_8 FILLER_26_1007 ();
 sg13g2_decap_8 FILLER_26_1014 ();
 sg13g2_decap_8 FILLER_26_1021 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_decap_4 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_fill_2 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_decap_4 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_94 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_4 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_446 ();
 sg13g2_decap_4 FILLER_27_465 ();
 sg13g2_fill_2 FILLER_27_474 ();
 sg13g2_decap_8 FILLER_27_519 ();
 sg13g2_decap_8 FILLER_27_526 ();
 sg13g2_decap_8 FILLER_27_533 ();
 sg13g2_decap_8 FILLER_27_540 ();
 sg13g2_fill_2 FILLER_27_547 ();
 sg13g2_fill_1 FILLER_27_549 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_fill_1 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_fill_2 FILLER_27_630 ();
 sg13g2_fill_1 FILLER_27_632 ();
 sg13g2_decap_8 FILLER_27_666 ();
 sg13g2_decap_4 FILLER_27_673 ();
 sg13g2_fill_1 FILLER_27_677 ();
 sg13g2_fill_1 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_730 ();
 sg13g2_decap_8 FILLER_27_737 ();
 sg13g2_decap_4 FILLER_27_744 ();
 sg13g2_fill_1 FILLER_27_748 ();
 sg13g2_fill_2 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_780 ();
 sg13g2_fill_2 FILLER_27_807 ();
 sg13g2_fill_1 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_853 ();
 sg13g2_decap_8 FILLER_27_860 ();
 sg13g2_decap_4 FILLER_27_867 ();
 sg13g2_fill_2 FILLER_27_871 ();
 sg13g2_fill_1 FILLER_27_885 ();
 sg13g2_fill_1 FILLER_27_895 ();
 sg13g2_fill_2 FILLER_27_901 ();
 sg13g2_fill_1 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_907 ();
 sg13g2_decap_8 FILLER_27_914 ();
 sg13g2_decap_8 FILLER_27_921 ();
 sg13g2_decap_8 FILLER_27_928 ();
 sg13g2_decap_8 FILLER_27_935 ();
 sg13g2_decap_8 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_decap_8 FILLER_27_956 ();
 sg13g2_decap_8 FILLER_27_963 ();
 sg13g2_decap_8 FILLER_27_970 ();
 sg13g2_decap_8 FILLER_27_977 ();
 sg13g2_decap_8 FILLER_27_984 ();
 sg13g2_decap_8 FILLER_27_991 ();
 sg13g2_decap_8 FILLER_27_998 ();
 sg13g2_decap_8 FILLER_27_1005 ();
 sg13g2_decap_8 FILLER_27_1012 ();
 sg13g2_decap_8 FILLER_27_1019 ();
 sg13g2_fill_2 FILLER_27_1026 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_2 FILLER_28_5 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_20 ();
 sg13g2_decap_8 FILLER_28_27 ();
 sg13g2_decap_8 FILLER_28_34 ();
 sg13g2_decap_8 FILLER_28_41 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_57 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_decap_8 FILLER_28_68 ();
 sg13g2_decap_4 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_decap_4 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_decap_8 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_decap_4 FILLER_28_320 ();
 sg13g2_decap_4 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_fill_2 FILLER_28_403 ();
 sg13g2_fill_1 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_28_436 ();
 sg13g2_fill_1 FILLER_28_443 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_decap_8 FILLER_28_471 ();
 sg13g2_decap_8 FILLER_28_478 ();
 sg13g2_decap_8 FILLER_28_489 ();
 sg13g2_decap_8 FILLER_28_496 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_fill_2 FILLER_28_517 ();
 sg13g2_fill_2 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_580 ();
 sg13g2_decap_4 FILLER_28_587 ();
 sg13g2_fill_2 FILLER_28_591 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_fill_2 FILLER_28_634 ();
 sg13g2_fill_1 FILLER_28_636 ();
 sg13g2_fill_2 FILLER_28_650 ();
 sg13g2_fill_1 FILLER_28_652 ();
 sg13g2_decap_4 FILLER_28_665 ();
 sg13g2_fill_1 FILLER_28_669 ();
 sg13g2_decap_4 FILLER_28_676 ();
 sg13g2_fill_2 FILLER_28_698 ();
 sg13g2_fill_1 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_4 FILLER_28_736 ();
 sg13g2_fill_1 FILLER_28_740 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_fill_2 FILLER_28_762 ();
 sg13g2_decap_4 FILLER_28_773 ();
 sg13g2_decap_4 FILLER_28_785 ();
 sg13g2_decap_8 FILLER_28_803 ();
 sg13g2_decap_4 FILLER_28_810 ();
 sg13g2_fill_2 FILLER_28_814 ();
 sg13g2_decap_4 FILLER_28_855 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_879 ();
 sg13g2_fill_1 FILLER_28_890 ();
 sg13g2_decap_8 FILLER_28_915 ();
 sg13g2_decap_8 FILLER_28_922 ();
 sg13g2_decap_8 FILLER_28_929 ();
 sg13g2_decap_8 FILLER_28_936 ();
 sg13g2_decap_8 FILLER_28_943 ();
 sg13g2_decap_8 FILLER_28_950 ();
 sg13g2_decap_8 FILLER_28_957 ();
 sg13g2_decap_8 FILLER_28_964 ();
 sg13g2_decap_8 FILLER_28_971 ();
 sg13g2_decap_8 FILLER_28_978 ();
 sg13g2_decap_8 FILLER_28_985 ();
 sg13g2_decap_8 FILLER_28_992 ();
 sg13g2_decap_8 FILLER_28_999 ();
 sg13g2_decap_8 FILLER_28_1006 ();
 sg13g2_decap_8 FILLER_28_1013 ();
 sg13g2_decap_8 FILLER_28_1020 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_2 FILLER_29_37 ();
 sg13g2_decap_8 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_decap_8 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_decap_4 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_158 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_decap_4 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_decap_4 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_261 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_4 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_372 ();
 sg13g2_decap_4 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_431 ();
 sg13g2_fill_2 FILLER_29_438 ();
 sg13g2_decap_8 FILLER_29_507 ();
 sg13g2_fill_1 FILLER_29_514 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_decap_8 FILLER_29_584 ();
 sg13g2_decap_8 FILLER_29_591 ();
 sg13g2_fill_2 FILLER_29_605 ();
 sg13g2_fill_1 FILLER_29_634 ();
 sg13g2_decap_4 FILLER_29_648 ();
 sg13g2_fill_2 FILLER_29_657 ();
 sg13g2_fill_1 FILLER_29_659 ();
 sg13g2_fill_2 FILLER_29_664 ();
 sg13g2_decap_4 FILLER_29_694 ();
 sg13g2_fill_2 FILLER_29_698 ();
 sg13g2_fill_2 FILLER_29_704 ();
 sg13g2_fill_1 FILLER_29_706 ();
 sg13g2_decap_4 FILLER_29_711 ();
 sg13g2_fill_1 FILLER_29_715 ();
 sg13g2_decap_8 FILLER_29_720 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_fill_1 FILLER_29_734 ();
 sg13g2_decap_4 FILLER_29_764 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_4 FILLER_29_783 ();
 sg13g2_fill_1 FILLER_29_787 ();
 sg13g2_decap_8 FILLER_29_813 ();
 sg13g2_decap_4 FILLER_29_820 ();
 sg13g2_fill_2 FILLER_29_824 ();
 sg13g2_fill_1 FILLER_29_838 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_fill_1 FILLER_29_865 ();
 sg13g2_decap_4 FILLER_29_883 ();
 sg13g2_fill_2 FILLER_29_887 ();
 sg13g2_fill_2 FILLER_29_895 ();
 sg13g2_decap_8 FILLER_29_916 ();
 sg13g2_decap_8 FILLER_29_923 ();
 sg13g2_decap_8 FILLER_29_930 ();
 sg13g2_decap_8 FILLER_29_937 ();
 sg13g2_decap_8 FILLER_29_944 ();
 sg13g2_decap_8 FILLER_29_951 ();
 sg13g2_decap_8 FILLER_29_958 ();
 sg13g2_decap_8 FILLER_29_965 ();
 sg13g2_decap_8 FILLER_29_972 ();
 sg13g2_decap_8 FILLER_29_979 ();
 sg13g2_decap_8 FILLER_29_986 ();
 sg13g2_decap_8 FILLER_29_993 ();
 sg13g2_decap_8 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1007 ();
 sg13g2_decap_8 FILLER_29_1014 ();
 sg13g2_decap_8 FILLER_29_1021 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_9 ();
 sg13g2_decap_4 FILLER_30_16 ();
 sg13g2_fill_2 FILLER_30_20 ();
 sg13g2_fill_2 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_94 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_decap_4 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_4 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_30_415 ();
 sg13g2_fill_2 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_424 ();
 sg13g2_decap_4 FILLER_30_464 ();
 sg13g2_fill_2 FILLER_30_468 ();
 sg13g2_decap_8 FILLER_30_484 ();
 sg13g2_decap_8 FILLER_30_491 ();
 sg13g2_fill_1 FILLER_30_498 ();
 sg13g2_decap_4 FILLER_30_503 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_fill_2 FILLER_30_518 ();
 sg13g2_fill_1 FILLER_30_524 ();
 sg13g2_fill_2 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_559 ();
 sg13g2_fill_2 FILLER_30_566 ();
 sg13g2_fill_1 FILLER_30_568 ();
 sg13g2_decap_8 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_580 ();
 sg13g2_decap_8 FILLER_30_587 ();
 sg13g2_decap_4 FILLER_30_594 ();
 sg13g2_fill_1 FILLER_30_598 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_4 FILLER_30_634 ();
 sg13g2_fill_2 FILLER_30_638 ();
 sg13g2_decap_4 FILLER_30_645 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_4 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_fill_1 FILLER_30_742 ();
 sg13g2_fill_1 FILLER_30_755 ();
 sg13g2_decap_4 FILLER_30_761 ();
 sg13g2_fill_1 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_fill_2 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_845 ();
 sg13g2_fill_2 FILLER_30_852 ();
 sg13g2_decap_8 FILLER_30_867 ();
 sg13g2_decap_4 FILLER_30_874 ();
 sg13g2_fill_1 FILLER_30_878 ();
 sg13g2_fill_1 FILLER_30_892 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_17 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_31 ();
 sg13g2_decap_8 FILLER_31_38 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_decap_4 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_decap_4 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_114 ();
 sg13g2_decap_8 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_138 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_decap_4 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_333 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_decap_4 FILLER_31_391 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_414 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_fill_2 FILLER_31_448 ();
 sg13g2_fill_1 FILLER_31_450 ();
 sg13g2_decap_8 FILLER_31_471 ();
 sg13g2_decap_4 FILLER_31_478 ();
 sg13g2_fill_2 FILLER_31_482 ();
 sg13g2_decap_4 FILLER_31_521 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_fill_2 FILLER_31_530 ();
 sg13g2_fill_1 FILLER_31_532 ();
 sg13g2_fill_2 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_fill_2 FILLER_31_592 ();
 sg13g2_fill_2 FILLER_31_602 ();
 sg13g2_decap_4 FILLER_31_608 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_fill_2 FILLER_31_651 ();
 sg13g2_fill_1 FILLER_31_653 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_fill_1 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_677 ();
 sg13g2_decap_4 FILLER_31_684 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_decap_8 FILLER_31_699 ();
 sg13g2_fill_2 FILLER_31_706 ();
 sg13g2_fill_1 FILLER_31_708 ();
 sg13g2_fill_2 FILLER_31_722 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_fill_2 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_fill_2 FILLER_31_769 ();
 sg13g2_fill_1 FILLER_31_771 ();
 sg13g2_decap_4 FILLER_31_788 ();
 sg13g2_fill_2 FILLER_31_792 ();
 sg13g2_decap_4 FILLER_31_815 ();
 sg13g2_fill_1 FILLER_31_847 ();
 sg13g2_fill_2 FILLER_31_851 ();
 sg13g2_fill_1 FILLER_31_853 ();
 sg13g2_fill_1 FILLER_31_880 ();
 sg13g2_decap_8 FILLER_31_900 ();
 sg13g2_decap_8 FILLER_31_907 ();
 sg13g2_decap_8 FILLER_31_914 ();
 sg13g2_decap_8 FILLER_31_921 ();
 sg13g2_decap_8 FILLER_31_928 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_8 FILLER_31_942 ();
 sg13g2_decap_8 FILLER_31_949 ();
 sg13g2_decap_8 FILLER_31_956 ();
 sg13g2_decap_8 FILLER_31_963 ();
 sg13g2_decap_8 FILLER_31_970 ();
 sg13g2_decap_8 FILLER_31_977 ();
 sg13g2_decap_8 FILLER_31_984 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_decap_8 FILLER_31_1005 ();
 sg13g2_decap_8 FILLER_31_1012 ();
 sg13g2_decap_8 FILLER_31_1019 ();
 sg13g2_fill_2 FILLER_31_1026 ();
 sg13g2_fill_1 FILLER_31_1028 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_decap_4 FILLER_32_345 ();
 sg13g2_decap_4 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_32_410 ();
 sg13g2_fill_2 FILLER_32_451 ();
 sg13g2_fill_1 FILLER_32_453 ();
 sg13g2_decap_8 FILLER_32_486 ();
 sg13g2_decap_4 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_497 ();
 sg13g2_fill_1 FILLER_32_507 ();
 sg13g2_decap_4 FILLER_32_525 ();
 sg13g2_fill_1 FILLER_32_529 ();
 sg13g2_fill_2 FILLER_32_557 ();
 sg13g2_fill_1 FILLER_32_559 ();
 sg13g2_decap_8 FILLER_32_568 ();
 sg13g2_decap_8 FILLER_32_575 ();
 sg13g2_fill_2 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_584 ();
 sg13g2_decap_8 FILLER_32_611 ();
 sg13g2_decap_8 FILLER_32_618 ();
 sg13g2_fill_2 FILLER_32_625 ();
 sg13g2_fill_1 FILLER_32_627 ();
 sg13g2_decap_8 FILLER_32_632 ();
 sg13g2_decap_8 FILLER_32_639 ();
 sg13g2_decap_8 FILLER_32_646 ();
 sg13g2_fill_1 FILLER_32_653 ();
 sg13g2_fill_1 FILLER_32_713 ();
 sg13g2_decap_8 FILLER_32_733 ();
 sg13g2_decap_8 FILLER_32_740 ();
 sg13g2_fill_2 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_764 ();
 sg13g2_fill_2 FILLER_32_771 ();
 sg13g2_decap_4 FILLER_32_783 ();
 sg13g2_fill_2 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_fill_2 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_fill_2 FILLER_32_857 ();
 sg13g2_fill_1 FILLER_32_859 ();
 sg13g2_decap_8 FILLER_32_874 ();
 sg13g2_fill_2 FILLER_32_881 ();
 sg13g2_fill_1 FILLER_32_883 ();
 sg13g2_decap_8 FILLER_32_922 ();
 sg13g2_decap_8 FILLER_32_929 ();
 sg13g2_decap_8 FILLER_32_936 ();
 sg13g2_decap_8 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_950 ();
 sg13g2_decap_8 FILLER_32_957 ();
 sg13g2_decap_8 FILLER_32_964 ();
 sg13g2_decap_8 FILLER_32_971 ();
 sg13g2_decap_8 FILLER_32_978 ();
 sg13g2_decap_8 FILLER_32_985 ();
 sg13g2_decap_8 FILLER_32_992 ();
 sg13g2_decap_8 FILLER_32_999 ();
 sg13g2_decap_8 FILLER_32_1006 ();
 sg13g2_decap_8 FILLER_32_1013 ();
 sg13g2_decap_4 FILLER_32_1020 ();
 sg13g2_fill_1 FILLER_32_1024 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_decap_4 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_51 ();
 sg13g2_fill_1 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_97 ();
 sg13g2_decap_8 FILLER_33_104 ();
 sg13g2_decap_8 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_decap_4 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_33_436 ();
 sg13g2_decap_8 FILLER_33_443 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_fill_1 FILLER_33_476 ();
 sg13g2_fill_1 FILLER_33_481 ();
 sg13g2_fill_1 FILLER_33_492 ();
 sg13g2_decap_8 FILLER_33_524 ();
 sg13g2_decap_8 FILLER_33_531 ();
 sg13g2_fill_2 FILLER_33_538 ();
 sg13g2_fill_1 FILLER_33_540 ();
 sg13g2_decap_8 FILLER_33_557 ();
 sg13g2_decap_8 FILLER_33_564 ();
 sg13g2_fill_2 FILLER_33_571 ();
 sg13g2_fill_1 FILLER_33_576 ();
 sg13g2_fill_1 FILLER_33_599 ();
 sg13g2_decap_8 FILLER_33_606 ();
 sg13g2_decap_8 FILLER_33_613 ();
 sg13g2_decap_8 FILLER_33_620 ();
 sg13g2_decap_4 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_635 ();
 sg13g2_decap_8 FILLER_33_642 ();
 sg13g2_decap_8 FILLER_33_649 ();
 sg13g2_decap_4 FILLER_33_656 ();
 sg13g2_decap_8 FILLER_33_664 ();
 sg13g2_decap_8 FILLER_33_671 ();
 sg13g2_decap_8 FILLER_33_678 ();
 sg13g2_fill_2 FILLER_33_685 ();
 sg13g2_decap_4 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_704 ();
 sg13g2_decap_4 FILLER_33_711 ();
 sg13g2_fill_2 FILLER_33_715 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_decap_8 FILLER_33_783 ();
 sg13g2_decap_4 FILLER_33_790 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_fill_2 FILLER_33_809 ();
 sg13g2_fill_1 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_fill_1 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_857 ();
 sg13g2_fill_2 FILLER_33_864 ();
 sg13g2_fill_1 FILLER_33_866 ();
 sg13g2_fill_2 FILLER_33_877 ();
 sg13g2_fill_1 FILLER_33_879 ();
 sg13g2_decap_8 FILLER_33_886 ();
 sg13g2_decap_4 FILLER_33_893 ();
 sg13g2_fill_2 FILLER_33_897 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_13 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_fill_2 FILLER_34_36 ();
 sg13g2_decap_8 FILLER_34_46 ();
 sg13g2_decap_4 FILLER_34_53 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_86 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_4 FILLER_34_177 ();
 sg13g2_fill_2 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_247 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_4 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_fill_1 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_decap_4 FILLER_34_440 ();
 sg13g2_decap_4 FILLER_34_476 ();
 sg13g2_fill_2 FILLER_34_490 ();
 sg13g2_fill_1 FILLER_34_492 ();
 sg13g2_decap_8 FILLER_34_520 ();
 sg13g2_decap_8 FILLER_34_527 ();
 sg13g2_decap_4 FILLER_34_534 ();
 sg13g2_fill_2 FILLER_34_546 ();
 sg13g2_fill_1 FILLER_34_548 ();
 sg13g2_fill_2 FILLER_34_564 ();
 sg13g2_fill_1 FILLER_34_566 ();
 sg13g2_fill_2 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_fill_2 FILLER_34_615 ();
 sg13g2_fill_1 FILLER_34_617 ();
 sg13g2_decap_8 FILLER_34_633 ();
 sg13g2_decap_8 FILLER_34_640 ();
 sg13g2_decap_4 FILLER_34_647 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_fill_2 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_4 FILLER_34_712 ();
 sg13g2_fill_2 FILLER_34_720 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_4 FILLER_34_747 ();
 sg13g2_fill_1 FILLER_34_751 ();
 sg13g2_fill_1 FILLER_34_761 ();
 sg13g2_fill_2 FILLER_34_816 ();
 sg13g2_fill_1 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_decap_8 FILLER_34_915 ();
 sg13g2_decap_8 FILLER_34_922 ();
 sg13g2_decap_8 FILLER_34_929 ();
 sg13g2_decap_8 FILLER_34_936 ();
 sg13g2_decap_8 FILLER_34_943 ();
 sg13g2_decap_8 FILLER_34_950 ();
 sg13g2_decap_8 FILLER_34_957 ();
 sg13g2_decap_8 FILLER_34_964 ();
 sg13g2_decap_8 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_decap_8 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1006 ();
 sg13g2_decap_8 FILLER_34_1013 ();
 sg13g2_decap_8 FILLER_34_1020 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_47 ();
 sg13g2_fill_2 FILLER_35_54 ();
 sg13g2_decap_4 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_4 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_decap_4 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_329 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_410 ();
 sg13g2_fill_1 FILLER_35_412 ();
 sg13g2_fill_2 FILLER_35_424 ();
 sg13g2_decap_8 FILLER_35_430 ();
 sg13g2_decap_8 FILLER_35_437 ();
 sg13g2_decap_4 FILLER_35_444 ();
 sg13g2_fill_1 FILLER_35_448 ();
 sg13g2_decap_4 FILLER_35_462 ();
 sg13g2_fill_2 FILLER_35_466 ();
 sg13g2_decap_8 FILLER_35_473 ();
 sg13g2_decap_8 FILLER_35_480 ();
 sg13g2_decap_8 FILLER_35_487 ();
 sg13g2_decap_4 FILLER_35_494 ();
 sg13g2_decap_4 FILLER_35_502 ();
 sg13g2_fill_1 FILLER_35_506 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_decap_8 FILLER_35_522 ();
 sg13g2_decap_4 FILLER_35_529 ();
 sg13g2_fill_2 FILLER_35_533 ();
 sg13g2_fill_1 FILLER_35_543 ();
 sg13g2_fill_2 FILLER_35_552 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_decap_4 FILLER_35_565 ();
 sg13g2_fill_2 FILLER_35_574 ();
 sg13g2_fill_1 FILLER_35_576 ();
 sg13g2_decap_8 FILLER_35_586 ();
 sg13g2_decap_4 FILLER_35_593 ();
 sg13g2_fill_2 FILLER_35_610 ();
 sg13g2_decap_4 FILLER_35_617 ();
 sg13g2_fill_1 FILLER_35_621 ();
 sg13g2_fill_1 FILLER_35_627 ();
 sg13g2_decap_4 FILLER_35_636 ();
 sg13g2_fill_2 FILLER_35_640 ();
 sg13g2_decap_8 FILLER_35_674 ();
 sg13g2_fill_1 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_fill_2 FILLER_35_794 ();
 sg13g2_fill_1 FILLER_35_823 ();
 sg13g2_decap_4 FILLER_35_828 ();
 sg13g2_fill_2 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_838 ();
 sg13g2_decap_8 FILLER_35_845 ();
 sg13g2_decap_4 FILLER_35_852 ();
 sg13g2_decap_8 FILLER_35_873 ();
 sg13g2_fill_1 FILLER_35_880 ();
 sg13g2_decap_4 FILLER_35_885 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_4 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_948 ();
 sg13g2_decap_8 FILLER_35_955 ();
 sg13g2_decap_8 FILLER_35_962 ();
 sg13g2_decap_8 FILLER_35_969 ();
 sg13g2_decap_8 FILLER_35_976 ();
 sg13g2_decap_8 FILLER_35_983 ();
 sg13g2_decap_8 FILLER_35_990 ();
 sg13g2_decap_8 FILLER_35_997 ();
 sg13g2_decap_8 FILLER_35_1004 ();
 sg13g2_decap_8 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1018 ();
 sg13g2_decap_4 FILLER_35_1025 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_decap_4 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_363 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_4 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_412 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_4 FILLER_36_448 ();
 sg13g2_fill_2 FILLER_36_452 ();
 sg13g2_decap_8 FILLER_36_468 ();
 sg13g2_decap_4 FILLER_36_475 ();
 sg13g2_fill_1 FILLER_36_493 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_decap_8 FILLER_36_528 ();
 sg13g2_fill_1 FILLER_36_535 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_decap_8 FILLER_36_555 ();
 sg13g2_fill_1 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_579 ();
 sg13g2_decap_8 FILLER_36_586 ();
 sg13g2_decap_4 FILLER_36_593 ();
 sg13g2_fill_1 FILLER_36_597 ();
 sg13g2_decap_8 FILLER_36_606 ();
 sg13g2_decap_8 FILLER_36_613 ();
 sg13g2_fill_1 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_4 FILLER_36_651 ();
 sg13g2_decap_4 FILLER_36_712 ();
 sg13g2_fill_1 FILLER_36_716 ();
 sg13g2_fill_1 FILLER_36_748 ();
 sg13g2_decap_8 FILLER_36_786 ();
 sg13g2_decap_8 FILLER_36_793 ();
 sg13g2_fill_1 FILLER_36_800 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_fill_2 FILLER_36_821 ();
 sg13g2_fill_1 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_4 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_878 ();
 sg13g2_decap_8 FILLER_36_885 ();
 sg13g2_fill_2 FILLER_36_892 ();
 sg13g2_decap_8 FILLER_36_898 ();
 sg13g2_fill_2 FILLER_36_905 ();
 sg13g2_decap_4 FILLER_36_920 ();
 sg13g2_fill_1 FILLER_36_924 ();
 sg13g2_fill_2 FILLER_36_937 ();
 sg13g2_fill_1 FILLER_36_939 ();
 sg13g2_fill_2 FILLER_36_947 ();
 sg13g2_decap_8 FILLER_36_962 ();
 sg13g2_decap_8 FILLER_36_969 ();
 sg13g2_decap_8 FILLER_36_976 ();
 sg13g2_decap_8 FILLER_36_983 ();
 sg13g2_decap_8 FILLER_36_990 ();
 sg13g2_decap_8 FILLER_36_997 ();
 sg13g2_decap_8 FILLER_36_1004 ();
 sg13g2_decap_8 FILLER_36_1011 ();
 sg13g2_decap_8 FILLER_36_1018 ();
 sg13g2_decap_4 FILLER_36_1025 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_12 ();
 sg13g2_fill_1 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_25 ();
 sg13g2_decap_8 FILLER_37_32 ();
 sg13g2_decap_4 FILLER_37_39 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_82 ();
 sg13g2_fill_1 FILLER_37_89 ();
 sg13g2_decap_4 FILLER_37_122 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_4 FILLER_37_161 ();
 sg13g2_decap_4 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_215 ();
 sg13g2_decap_4 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_decap_4 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_396 ();
 sg13g2_fill_1 FILLER_37_398 ();
 sg13g2_fill_1 FILLER_37_475 ();
 sg13g2_decap_8 FILLER_37_491 ();
 sg13g2_fill_2 FILLER_37_498 ();
 sg13g2_decap_4 FILLER_37_504 ();
 sg13g2_fill_1 FILLER_37_513 ();
 sg13g2_fill_2 FILLER_37_527 ();
 sg13g2_fill_1 FILLER_37_529 ();
 sg13g2_decap_4 FILLER_37_573 ();
 sg13g2_fill_1 FILLER_37_577 ();
 sg13g2_decap_8 FILLER_37_586 ();
 sg13g2_fill_2 FILLER_37_614 ();
 sg13g2_decap_8 FILLER_37_641 ();
 sg13g2_fill_2 FILLER_37_648 ();
 sg13g2_fill_1 FILLER_37_650 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_fill_1 FILLER_37_706 ();
 sg13g2_decap_4 FILLER_37_726 ();
 sg13g2_decap_4 FILLER_37_753 ();
 sg13g2_fill_1 FILLER_37_757 ();
 sg13g2_decap_8 FILLER_37_768 ();
 sg13g2_decap_8 FILLER_37_775 ();
 sg13g2_fill_1 FILLER_37_782 ();
 sg13g2_fill_1 FILLER_37_820 ();
 sg13g2_decap_4 FILLER_37_858 ();
 sg13g2_fill_2 FILLER_37_862 ();
 sg13g2_decap_8 FILLER_37_897 ();
 sg13g2_fill_2 FILLER_37_904 ();
 sg13g2_fill_1 FILLER_37_906 ();
 sg13g2_decap_8 FILLER_37_922 ();
 sg13g2_decap_4 FILLER_37_929 ();
 sg13g2_decap_4 FILLER_37_960 ();
 sg13g2_decap_8 FILLER_37_972 ();
 sg13g2_decap_8 FILLER_37_979 ();
 sg13g2_decap_8 FILLER_37_986 ();
 sg13g2_decap_8 FILLER_37_993 ();
 sg13g2_decap_8 FILLER_37_1000 ();
 sg13g2_decap_8 FILLER_37_1007 ();
 sg13g2_decap_8 FILLER_37_1014 ();
 sg13g2_decap_8 FILLER_37_1021 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_decap_4 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_fill_2 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_58 ();
 sg13g2_decap_8 FILLER_38_67 ();
 sg13g2_decap_8 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_81 ();
 sg13g2_decap_8 FILLER_38_88 ();
 sg13g2_decap_4 FILLER_38_99 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_decap_8 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_115 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_141 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_decap_4 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_405 ();
 sg13g2_fill_1 FILLER_38_407 ();
 sg13g2_decap_4 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_426 ();
 sg13g2_fill_2 FILLER_38_433 ();
 sg13g2_fill_1 FILLER_38_445 ();
 sg13g2_decap_4 FILLER_38_450 ();
 sg13g2_fill_2 FILLER_38_459 ();
 sg13g2_fill_1 FILLER_38_461 ();
 sg13g2_decap_4 FILLER_38_480 ();
 sg13g2_fill_2 FILLER_38_484 ();
 sg13g2_decap_4 FILLER_38_496 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_decap_4 FILLER_38_586 ();
 sg13g2_fill_1 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_616 ();
 sg13g2_fill_1 FILLER_38_618 ();
 sg13g2_decap_8 FILLER_38_633 ();
 sg13g2_decap_8 FILLER_38_640 ();
 sg13g2_decap_8 FILLER_38_647 ();
 sg13g2_decap_4 FILLER_38_654 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_704 ();
 sg13g2_fill_2 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_846 ();
 sg13g2_fill_2 FILLER_38_853 ();
 sg13g2_fill_1 FILLER_38_855 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_38_867 ();
 sg13g2_decap_8 FILLER_38_874 ();
 sg13g2_decap_8 FILLER_38_881 ();
 sg13g2_fill_2 FILLER_38_888 ();
 sg13g2_fill_1 FILLER_38_890 ();
 sg13g2_decap_4 FILLER_38_901 ();
 sg13g2_fill_1 FILLER_38_905 ();
 sg13g2_fill_1 FILLER_38_923 ();
 sg13g2_fill_2 FILLER_38_938 ();
 sg13g2_decap_4 FILLER_38_958 ();
 sg13g2_decap_8 FILLER_38_972 ();
 sg13g2_decap_8 FILLER_38_979 ();
 sg13g2_decap_8 FILLER_38_986 ();
 sg13g2_decap_8 FILLER_38_993 ();
 sg13g2_decap_8 FILLER_38_1000 ();
 sg13g2_decap_8 FILLER_38_1007 ();
 sg13g2_decap_8 FILLER_38_1014 ();
 sg13g2_decap_8 FILLER_38_1021 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_12 ();
 sg13g2_decap_8 FILLER_39_20 ();
 sg13g2_decap_8 FILLER_39_27 ();
 sg13g2_decap_4 FILLER_39_34 ();
 sg13g2_decap_8 FILLER_39_48 ();
 sg13g2_fill_2 FILLER_39_55 ();
 sg13g2_fill_1 FILLER_39_57 ();
 sg13g2_fill_1 FILLER_39_62 ();
 sg13g2_fill_1 FILLER_39_76 ();
 sg13g2_decap_8 FILLER_39_102 ();
 sg13g2_fill_2 FILLER_39_113 ();
 sg13g2_decap_4 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_decap_4 FILLER_39_187 ();
 sg13g2_decap_8 FILLER_39_218 ();
 sg13g2_fill_2 FILLER_39_225 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_232 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_277 ();
 sg13g2_decap_4 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_300 ();
 sg13g2_decap_8 FILLER_39_309 ();
 sg13g2_decap_8 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_323 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_decap_4 FILLER_39_341 ();
 sg13g2_decap_8 FILLER_39_349 ();
 sg13g2_decap_8 FILLER_39_356 ();
 sg13g2_decap_8 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_1 FILLER_39_391 ();
 sg13g2_decap_4 FILLER_39_431 ();
 sg13g2_fill_1 FILLER_39_462 ();
 sg13g2_decap_4 FILLER_39_500 ();
 sg13g2_fill_1 FILLER_39_504 ();
 sg13g2_decap_4 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_517 ();
 sg13g2_decap_8 FILLER_39_524 ();
 sg13g2_decap_8 FILLER_39_531 ();
 sg13g2_fill_2 FILLER_39_538 ();
 sg13g2_decap_4 FILLER_39_560 ();
 sg13g2_fill_2 FILLER_39_564 ();
 sg13g2_decap_8 FILLER_39_585 ();
 sg13g2_fill_2 FILLER_39_592 ();
 sg13g2_fill_1 FILLER_39_594 ();
 sg13g2_decap_8 FILLER_39_605 ();
 sg13g2_fill_2 FILLER_39_618 ();
 sg13g2_fill_1 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_645 ();
 sg13g2_decap_8 FILLER_39_652 ();
 sg13g2_decap_8 FILLER_39_659 ();
 sg13g2_decap_4 FILLER_39_666 ();
 sg13g2_fill_1 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_706 ();
 sg13g2_fill_1 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_fill_1 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_750 ();
 sg13g2_decap_4 FILLER_39_757 ();
 sg13g2_fill_2 FILLER_39_761 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_fill_1 FILLER_39_784 ();
 sg13g2_decap_4 FILLER_39_804 ();
 sg13g2_fill_1 FILLER_39_808 ();
 sg13g2_decap_8 FILLER_39_838 ();
 sg13g2_decap_4 FILLER_39_845 ();
 sg13g2_fill_1 FILLER_39_849 ();
 sg13g2_fill_2 FILLER_39_855 ();
 sg13g2_fill_1 FILLER_39_857 ();
 sg13g2_decap_8 FILLER_39_883 ();
 sg13g2_fill_2 FILLER_39_890 ();
 sg13g2_fill_1 FILLER_39_892 ();
 sg13g2_fill_2 FILLER_39_901 ();
 sg13g2_fill_1 FILLER_39_903 ();
 sg13g2_fill_2 FILLER_39_912 ();
 sg13g2_decap_8 FILLER_39_932 ();
 sg13g2_decap_8 FILLER_39_939 ();
 sg13g2_fill_2 FILLER_39_946 ();
 sg13g2_fill_1 FILLER_39_964 ();
 sg13g2_decap_8 FILLER_39_976 ();
 sg13g2_decap_8 FILLER_39_983 ();
 sg13g2_decap_8 FILLER_39_990 ();
 sg13g2_decap_8 FILLER_39_997 ();
 sg13g2_decap_8 FILLER_39_1004 ();
 sg13g2_decap_8 FILLER_39_1011 ();
 sg13g2_decap_8 FILLER_39_1018 ();
 sg13g2_decap_4 FILLER_39_1025 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_2 FILLER_40_40 ();
 sg13g2_fill_1 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_92 ();
 sg13g2_decap_8 FILLER_40_145 ();
 sg13g2_decap_4 FILLER_40_152 ();
 sg13g2_fill_2 FILLER_40_156 ();
 sg13g2_decap_4 FILLER_40_162 ();
 sg13g2_fill_2 FILLER_40_166 ();
 sg13g2_decap_8 FILLER_40_176 ();
 sg13g2_decap_8 FILLER_40_183 ();
 sg13g2_fill_2 FILLER_40_190 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_fill_2 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_259 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_313 ();
 sg13g2_decap_8 FILLER_40_320 ();
 sg13g2_decap_8 FILLER_40_367 ();
 sg13g2_decap_4 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_396 ();
 sg13g2_fill_2 FILLER_40_414 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_fill_2 FILLER_40_438 ();
 sg13g2_decap_8 FILLER_40_444 ();
 sg13g2_decap_8 FILLER_40_451 ();
 sg13g2_decap_8 FILLER_40_458 ();
 sg13g2_decap_8 FILLER_40_465 ();
 sg13g2_fill_2 FILLER_40_472 ();
 sg13g2_decap_8 FILLER_40_482 ();
 sg13g2_decap_8 FILLER_40_489 ();
 sg13g2_decap_8 FILLER_40_496 ();
 sg13g2_fill_2 FILLER_40_503 ();
 sg13g2_fill_1 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_4 FILLER_40_546 ();
 sg13g2_fill_2 FILLER_40_575 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_fill_1 FILLER_40_602 ();
 sg13g2_decap_4 FILLER_40_607 ();
 sg13g2_fill_2 FILLER_40_611 ();
 sg13g2_fill_2 FILLER_40_633 ();
 sg13g2_fill_1 FILLER_40_635 ();
 sg13g2_fill_1 FILLER_40_701 ();
 sg13g2_fill_2 FILLER_40_711 ();
 sg13g2_fill_1 FILLER_40_713 ();
 sg13g2_fill_2 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_792 ();
 sg13g2_fill_1 FILLER_40_799 ();
 sg13g2_decap_4 FILLER_40_831 ();
 sg13g2_fill_1 FILLER_40_835 ();
 sg13g2_decap_4 FILLER_40_883 ();
 sg13g2_fill_2 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_decap_4 FILLER_40_901 ();
 sg13g2_fill_2 FILLER_40_905 ();
 sg13g2_fill_1 FILLER_40_928 ();
 sg13g2_fill_2 FILLER_40_932 ();
 sg13g2_decap_8 FILLER_40_978 ();
 sg13g2_decap_8 FILLER_40_985 ();
 sg13g2_decap_8 FILLER_40_992 ();
 sg13g2_decap_8 FILLER_40_999 ();
 sg13g2_decap_8 FILLER_40_1006 ();
 sg13g2_decap_8 FILLER_40_1013 ();
 sg13g2_decap_8 FILLER_40_1020 ();
 sg13g2_fill_2 FILLER_40_1027 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_36 ();
 sg13g2_decap_8 FILLER_41_48 ();
 sg13g2_decap_8 FILLER_41_55 ();
 sg13g2_decap_4 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_87 ();
 sg13g2_decap_4 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_98 ();
 sg13g2_decap_4 FILLER_41_103 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_decap_4 FILLER_41_125 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_1 FILLER_41_151 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_decap_8 FILLER_41_243 ();
 sg13g2_decap_8 FILLER_41_250 ();
 sg13g2_fill_2 FILLER_41_257 ();
 sg13g2_fill_1 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_fill_2 FILLER_41_273 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_decap_8 FILLER_41_295 ();
 sg13g2_decap_4 FILLER_41_302 ();
 sg13g2_decap_4 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_324 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_fill_1 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_decap_8 FILLER_41_408 ();
 sg13g2_decap_4 FILLER_41_415 ();
 sg13g2_decap_4 FILLER_41_446 ();
 sg13g2_fill_1 FILLER_41_464 ();
 sg13g2_fill_1 FILLER_41_475 ();
 sg13g2_decap_4 FILLER_41_486 ();
 sg13g2_decap_4 FILLER_41_500 ();
 sg13g2_fill_1 FILLER_41_504 ();
 sg13g2_fill_2 FILLER_41_532 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_fill_2 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_fill_2 FILLER_41_569 ();
 sg13g2_fill_1 FILLER_41_571 ();
 sg13g2_decap_8 FILLER_41_600 ();
 sg13g2_decap_8 FILLER_41_607 ();
 sg13g2_decap_4 FILLER_41_624 ();
 sg13g2_fill_2 FILLER_41_628 ();
 sg13g2_fill_2 FILLER_41_662 ();
 sg13g2_decap_8 FILLER_41_709 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_fill_2 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_823 ();
 sg13g2_decap_8 FILLER_41_834 ();
 sg13g2_decap_8 FILLER_41_841 ();
 sg13g2_fill_2 FILLER_41_848 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_fill_2 FILLER_41_862 ();
 sg13g2_fill_1 FILLER_41_864 ();
 sg13g2_decap_4 FILLER_41_911 ();
 sg13g2_fill_2 FILLER_41_915 ();
 sg13g2_fill_2 FILLER_41_922 ();
 sg13g2_decap_4 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_972 ();
 sg13g2_decap_8 FILLER_41_979 ();
 sg13g2_decap_8 FILLER_41_986 ();
 sg13g2_decap_8 FILLER_41_993 ();
 sg13g2_decap_8 FILLER_41_1000 ();
 sg13g2_decap_8 FILLER_41_1007 ();
 sg13g2_decap_8 FILLER_41_1014 ();
 sg13g2_decap_8 FILLER_41_1021 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_11 ();
 sg13g2_decap_8 FILLER_42_29 ();
 sg13g2_decap_4 FILLER_42_36 ();
 sg13g2_fill_1 FILLER_42_40 ();
 sg13g2_decap_4 FILLER_42_46 ();
 sg13g2_fill_2 FILLER_42_77 ();
 sg13g2_fill_1 FILLER_42_79 ();
 sg13g2_decap_8 FILLER_42_121 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_fill_1 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_fill_1 FILLER_42_229 ();
 sg13g2_decap_8 FILLER_42_234 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_255 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_4 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_decap_4 FILLER_42_300 ();
 sg13g2_decap_4 FILLER_42_331 ();
 sg13g2_decap_8 FILLER_42_340 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_decap_8 FILLER_42_354 ();
 sg13g2_fill_2 FILLER_42_361 ();
 sg13g2_fill_1 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_400 ();
 sg13g2_decap_4 FILLER_42_407 ();
 sg13g2_decap_4 FILLER_42_421 ();
 sg13g2_fill_1 FILLER_42_425 ();
 sg13g2_decap_8 FILLER_42_457 ();
 sg13g2_decap_4 FILLER_42_464 ();
 sg13g2_fill_2 FILLER_42_468 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_4 FILLER_42_504 ();
 sg13g2_fill_2 FILLER_42_508 ();
 sg13g2_fill_2 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_516 ();
 sg13g2_decap_4 FILLER_42_521 ();
 sg13g2_fill_1 FILLER_42_525 ();
 sg13g2_fill_1 FILLER_42_530 ();
 sg13g2_fill_1 FILLER_42_548 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_decap_8 FILLER_42_559 ();
 sg13g2_decap_8 FILLER_42_648 ();
 sg13g2_fill_2 FILLER_42_655 ();
 sg13g2_decap_4 FILLER_42_703 ();
 sg13g2_fill_1 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_730 ();
 sg13g2_fill_1 FILLER_42_737 ();
 sg13g2_decap_8 FILLER_42_751 ();
 sg13g2_decap_8 FILLER_42_758 ();
 sg13g2_fill_2 FILLER_42_765 ();
 sg13g2_fill_1 FILLER_42_767 ();
 sg13g2_fill_1 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_4 FILLER_42_867 ();
 sg13g2_fill_1 FILLER_42_871 ();
 sg13g2_decap_8 FILLER_42_885 ();
 sg13g2_decap_8 FILLER_42_892 ();
 sg13g2_decap_4 FILLER_42_899 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_966 ();
 sg13g2_decap_8 FILLER_42_973 ();
 sg13g2_decap_8 FILLER_42_980 ();
 sg13g2_decap_8 FILLER_42_987 ();
 sg13g2_decap_8 FILLER_42_994 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_44 ();
 sg13g2_decap_4 FILLER_43_50 ();
 sg13g2_fill_1 FILLER_43_54 ();
 sg13g2_fill_2 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_69 ();
 sg13g2_decap_4 FILLER_43_90 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_120 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_decap_4 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_194 ();
 sg13g2_decap_4 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_205 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_4 FILLER_43_256 ();
 sg13g2_fill_2 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_266 ();
 sg13g2_fill_1 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_fill_2 FILLER_43_287 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_fill_2 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_decap_4 FILLER_43_324 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_decap_8 FILLER_43_335 ();
 sg13g2_decap_8 FILLER_43_342 ();
 sg13g2_decap_4 FILLER_43_349 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_decap_4 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_384 ();
 sg13g2_fill_1 FILLER_43_389 ();
 sg13g2_fill_2 FILLER_43_422 ();
 sg13g2_decap_8 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_43_435 ();
 sg13g2_fill_2 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_442 ();
 sg13g2_decap_8 FILLER_43_447 ();
 sg13g2_fill_2 FILLER_43_454 ();
 sg13g2_decap_8 FILLER_43_465 ();
 sg13g2_fill_2 FILLER_43_472 ();
 sg13g2_fill_1 FILLER_43_474 ();
 sg13g2_fill_2 FILLER_43_479 ();
 sg13g2_fill_2 FILLER_43_485 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_decap_4 FILLER_43_492 ();
 sg13g2_fill_2 FILLER_43_496 ();
 sg13g2_fill_2 FILLER_43_511 ();
 sg13g2_fill_1 FILLER_43_513 ();
 sg13g2_decap_8 FILLER_43_541 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_8 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_fill_2 FILLER_43_569 ();
 sg13g2_decap_8 FILLER_43_575 ();
 sg13g2_decap_8 FILLER_43_582 ();
 sg13g2_decap_4 FILLER_43_594 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_4 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_4 FILLER_43_635 ();
 sg13g2_fill_1 FILLER_43_639 ();
 sg13g2_fill_2 FILLER_43_644 ();
 sg13g2_fill_2 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_fill_2 FILLER_43_773 ();
 sg13g2_fill_1 FILLER_43_775 ();
 sg13g2_decap_4 FILLER_43_789 ();
 sg13g2_fill_1 FILLER_43_819 ();
 sg13g2_decap_4 FILLER_43_901 ();
 sg13g2_fill_1 FILLER_43_905 ();
 sg13g2_decap_8 FILLER_43_934 ();
 sg13g2_decap_8 FILLER_43_941 ();
 sg13g2_decap_8 FILLER_43_948 ();
 sg13g2_decap_8 FILLER_43_955 ();
 sg13g2_decap_8 FILLER_43_962 ();
 sg13g2_decap_8 FILLER_43_969 ();
 sg13g2_decap_8 FILLER_43_976 ();
 sg13g2_decap_8 FILLER_43_983 ();
 sg13g2_decap_8 FILLER_43_990 ();
 sg13g2_decap_8 FILLER_43_997 ();
 sg13g2_decap_8 FILLER_43_1004 ();
 sg13g2_decap_8 FILLER_43_1011 ();
 sg13g2_decap_8 FILLER_43_1018 ();
 sg13g2_decap_4 FILLER_43_1025 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_4 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_110 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_decap_4 FILLER_44_144 ();
 sg13g2_fill_2 FILLER_44_148 ();
 sg13g2_decap_4 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_198 ();
 sg13g2_decap_4 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_231 ();
 sg13g2_fill_1 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_245 ();
 sg13g2_decap_4 FILLER_44_270 ();
 sg13g2_fill_1 FILLER_44_274 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_fill_2 FILLER_44_362 ();
 sg13g2_decap_4 FILLER_44_391 ();
 sg13g2_fill_2 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_421 ();
 sg13g2_decap_4 FILLER_44_428 ();
 sg13g2_fill_1 FILLER_44_432 ();
 sg13g2_fill_2 FILLER_44_437 ();
 sg13g2_fill_1 FILLER_44_439 ();
 sg13g2_decap_4 FILLER_44_444 ();
 sg13g2_fill_1 FILLER_44_448 ();
 sg13g2_decap_4 FILLER_44_470 ();
 sg13g2_fill_1 FILLER_44_474 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_fill_2 FILLER_44_494 ();
 sg13g2_fill_2 FILLER_44_516 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_decap_4 FILLER_44_554 ();
 sg13g2_fill_2 FILLER_44_558 ();
 sg13g2_decap_4 FILLER_44_587 ();
 sg13g2_fill_1 FILLER_44_591 ();
 sg13g2_fill_1 FILLER_44_623 ();
 sg13g2_fill_1 FILLER_44_651 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_decap_8 FILLER_44_722 ();
 sg13g2_fill_2 FILLER_44_729 ();
 sg13g2_fill_1 FILLER_44_741 ();
 sg13g2_decap_4 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_773 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_4 FILLER_44_858 ();
 sg13g2_fill_1 FILLER_44_862 ();
 sg13g2_decap_8 FILLER_44_890 ();
 sg13g2_decap_8 FILLER_44_897 ();
 sg13g2_fill_2 FILLER_44_904 ();
 sg13g2_fill_1 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_915 ();
 sg13g2_decap_8 FILLER_44_922 ();
 sg13g2_decap_8 FILLER_44_929 ();
 sg13g2_decap_8 FILLER_44_936 ();
 sg13g2_decap_8 FILLER_44_943 ();
 sg13g2_decap_8 FILLER_44_950 ();
 sg13g2_decap_8 FILLER_44_957 ();
 sg13g2_decap_8 FILLER_44_964 ();
 sg13g2_decap_8 FILLER_44_971 ();
 sg13g2_decap_8 FILLER_44_978 ();
 sg13g2_decap_8 FILLER_44_985 ();
 sg13g2_decap_8 FILLER_44_992 ();
 sg13g2_decap_8 FILLER_44_999 ();
 sg13g2_decap_8 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1013 ();
 sg13g2_decap_8 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_25 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_fill_1 FILLER_45_34 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_60 ();
 sg13g2_decap_8 FILLER_45_66 ();
 sg13g2_fill_2 FILLER_45_73 ();
 sg13g2_fill_1 FILLER_45_75 ();
 sg13g2_fill_2 FILLER_45_86 ();
 sg13g2_decap_8 FILLER_45_92 ();
 sg13g2_decap_4 FILLER_45_99 ();
 sg13g2_decap_8 FILLER_45_142 ();
 sg13g2_decap_8 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_156 ();
 sg13g2_decap_4 FILLER_45_163 ();
 sg13g2_fill_2 FILLER_45_167 ();
 sg13g2_fill_2 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_175 ();
 sg13g2_decap_4 FILLER_45_180 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_8 FILLER_45_235 ();
 sg13g2_fill_2 FILLER_45_273 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_fill_1 FILLER_45_314 ();
 sg13g2_fill_2 FILLER_45_362 ();
 sg13g2_decap_8 FILLER_45_391 ();
 sg13g2_decap_4 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_407 ();
 sg13g2_fill_2 FILLER_45_470 ();
 sg13g2_fill_2 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_498 ();
 sg13g2_fill_2 FILLER_45_526 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_decap_8 FILLER_45_537 ();
 sg13g2_decap_8 FILLER_45_544 ();
 sg13g2_decap_8 FILLER_45_551 ();
 sg13g2_decap_8 FILLER_45_558 ();
 sg13g2_decap_8 FILLER_45_569 ();
 sg13g2_decap_8 FILLER_45_603 ();
 sg13g2_fill_1 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_615 ();
 sg13g2_fill_1 FILLER_45_617 ();
 sg13g2_decap_8 FILLER_45_631 ();
 sg13g2_decap_8 FILLER_45_638 ();
 sg13g2_decap_4 FILLER_45_645 ();
 sg13g2_fill_1 FILLER_45_649 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_fill_2 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_672 ();
 sg13g2_fill_2 FILLER_45_709 ();
 sg13g2_fill_1 FILLER_45_711 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_fill_1 FILLER_45_746 ();
 sg13g2_decap_4 FILLER_45_751 ();
 sg13g2_fill_2 FILLER_45_755 ();
 sg13g2_decap_4 FILLER_45_816 ();
 sg13g2_fill_2 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_fill_2 FILLER_45_865 ();
 sg13g2_fill_1 FILLER_45_867 ();
 sg13g2_decap_8 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_886 ();
 sg13g2_decap_8 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_914 ();
 sg13g2_decap_8 FILLER_45_921 ();
 sg13g2_decap_8 FILLER_45_928 ();
 sg13g2_decap_8 FILLER_45_935 ();
 sg13g2_decap_8 FILLER_45_942 ();
 sg13g2_decap_8 FILLER_45_949 ();
 sg13g2_decap_8 FILLER_45_956 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_8 FILLER_45_970 ();
 sg13g2_decap_8 FILLER_45_977 ();
 sg13g2_decap_8 FILLER_45_984 ();
 sg13g2_decap_8 FILLER_45_991 ();
 sg13g2_decap_8 FILLER_45_998 ();
 sg13g2_decap_8 FILLER_45_1005 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_4 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1023 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_25 ();
 sg13g2_decap_8 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_88 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_2 FILLER_46_172 ();
 sg13g2_fill_1 FILLER_46_174 ();
 sg13g2_decap_4 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_233 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_4 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_280 ();
 sg13g2_decap_4 FILLER_46_286 ();
 sg13g2_fill_2 FILLER_46_294 ();
 sg13g2_fill_1 FILLER_46_296 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_4 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_312 ();
 sg13g2_decap_8 FILLER_46_330 ();
 sg13g2_decap_4 FILLER_46_337 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_decap_4 FILLER_46_351 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_fill_2 FILLER_46_366 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_decap_4 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_4 FILLER_46_390 ();
 sg13g2_fill_2 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_422 ();
 sg13g2_decap_8 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_46_436 ();
 sg13g2_fill_2 FILLER_46_443 ();
 sg13g2_fill_1 FILLER_46_445 ();
 sg13g2_decap_8 FILLER_46_450 ();
 sg13g2_decap_4 FILLER_46_467 ();
 sg13g2_fill_1 FILLER_46_475 ();
 sg13g2_decap_8 FILLER_46_480 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_decap_4 FILLER_46_494 ();
 sg13g2_decap_8 FILLER_46_512 ();
 sg13g2_fill_2 FILLER_46_519 ();
 sg13g2_fill_1 FILLER_46_521 ();
 sg13g2_decap_8 FILLER_46_549 ();
 sg13g2_decap_8 FILLER_46_556 ();
 sg13g2_decap_8 FILLER_46_563 ();
 sg13g2_decap_8 FILLER_46_570 ();
 sg13g2_decap_8 FILLER_46_594 ();
 sg13g2_fill_2 FILLER_46_601 ();
 sg13g2_fill_2 FILLER_46_684 ();
 sg13g2_fill_1 FILLER_46_686 ();
 sg13g2_fill_1 FILLER_46_706 ();
 sg13g2_decap_8 FILLER_46_743 ();
 sg13g2_decap_4 FILLER_46_750 ();
 sg13g2_decap_4 FILLER_46_767 ();
 sg13g2_fill_1 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_decap_8 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_46_867 ();
 sg13g2_decap_8 FILLER_46_874 ();
 sg13g2_decap_8 FILLER_46_881 ();
 sg13g2_decap_8 FILLER_46_888 ();
 sg13g2_decap_8 FILLER_46_895 ();
 sg13g2_decap_8 FILLER_46_902 ();
 sg13g2_decap_8 FILLER_46_909 ();
 sg13g2_decap_8 FILLER_46_916 ();
 sg13g2_decap_8 FILLER_46_923 ();
 sg13g2_decap_8 FILLER_46_930 ();
 sg13g2_decap_8 FILLER_46_937 ();
 sg13g2_decap_8 FILLER_46_944 ();
 sg13g2_decap_8 FILLER_46_951 ();
 sg13g2_decap_8 FILLER_46_958 ();
 sg13g2_decap_8 FILLER_46_965 ();
 sg13g2_decap_8 FILLER_46_972 ();
 sg13g2_decap_8 FILLER_46_979 ();
 sg13g2_decap_8 FILLER_46_986 ();
 sg13g2_decap_8 FILLER_46_993 ();
 sg13g2_decap_8 FILLER_46_1000 ();
 sg13g2_decap_8 FILLER_46_1007 ();
 sg13g2_decap_8 FILLER_46_1014 ();
 sg13g2_decap_8 FILLER_46_1021 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_4 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_32 ();
 sg13g2_decap_8 FILLER_47_37 ();
 sg13g2_decap_8 FILLER_47_44 ();
 sg13g2_decap_8 FILLER_47_51 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_114 ();
 sg13g2_decap_4 FILLER_47_121 ();
 sg13g2_fill_2 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_141 ();
 sg13g2_decap_4 FILLER_47_148 ();
 sg13g2_decap_4 FILLER_47_206 ();
 sg13g2_fill_2 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_256 ();
 sg13g2_decap_4 FILLER_47_274 ();
 sg13g2_fill_2 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_290 ();
 sg13g2_decap_4 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_decap_4 FILLER_47_314 ();
 sg13g2_decap_4 FILLER_47_331 ();
 sg13g2_fill_1 FILLER_47_335 ();
 sg13g2_fill_2 FILLER_47_378 ();
 sg13g2_fill_1 FILLER_47_380 ();
 sg13g2_decap_4 FILLER_47_394 ();
 sg13g2_fill_2 FILLER_47_398 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_fill_2 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_440 ();
 sg13g2_decap_8 FILLER_47_446 ();
 sg13g2_decap_4 FILLER_47_453 ();
 sg13g2_fill_1 FILLER_47_457 ();
 sg13g2_fill_2 FILLER_47_525 ();
 sg13g2_fill_1 FILLER_47_531 ();
 sg13g2_decap_8 FILLER_47_536 ();
 sg13g2_decap_8 FILLER_47_543 ();
 sg13g2_decap_8 FILLER_47_550 ();
 sg13g2_decap_8 FILLER_47_557 ();
 sg13g2_decap_8 FILLER_47_564 ();
 sg13g2_decap_4 FILLER_47_571 ();
 sg13g2_fill_2 FILLER_47_575 ();
 sg13g2_decap_8 FILLER_47_582 ();
 sg13g2_decap_8 FILLER_47_589 ();
 sg13g2_fill_2 FILLER_47_596 ();
 sg13g2_fill_1 FILLER_47_598 ();
 sg13g2_decap_8 FILLER_47_613 ();
 sg13g2_decap_8 FILLER_47_620 ();
 sg13g2_fill_2 FILLER_47_627 ();
 sg13g2_decap_8 FILLER_47_643 ();
 sg13g2_decap_4 FILLER_47_650 ();
 sg13g2_fill_2 FILLER_47_654 ();
 sg13g2_fill_2 FILLER_47_683 ();
 sg13g2_decap_4 FILLER_47_742 ();
 sg13g2_fill_2 FILLER_47_746 ();
 sg13g2_decap_4 FILLER_47_775 ();
 sg13g2_decap_8 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_813 ();
 sg13g2_decap_8 FILLER_47_820 ();
 sg13g2_fill_1 FILLER_47_827 ();
 sg13g2_fill_2 FILLER_47_831 ();
 sg13g2_fill_1 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_decap_8 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_871 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_8 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_983 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_96 ();
 sg13g2_decap_8 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_decap_4 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_decap_8 FILLER_48_195 ();
 sg13g2_decap_8 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_209 ();
 sg13g2_decap_8 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_4 FILLER_48_401 ();
 sg13g2_decap_8 FILLER_48_409 ();
 sg13g2_fill_2 FILLER_48_416 ();
 sg13g2_fill_1 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_524 ();
 sg13g2_decap_8 FILLER_48_531 ();
 sg13g2_decap_8 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_545 ();
 sg13g2_decap_8 FILLER_48_552 ();
 sg13g2_decap_8 FILLER_48_559 ();
 sg13g2_decap_8 FILLER_48_566 ();
 sg13g2_decap_4 FILLER_48_573 ();
 sg13g2_fill_2 FILLER_48_577 ();
 sg13g2_fill_1 FILLER_48_606 ();
 sg13g2_decap_4 FILLER_48_634 ();
 sg13g2_fill_1 FILLER_48_638 ();
 sg13g2_decap_8 FILLER_48_666 ();
 sg13g2_fill_1 FILLER_48_709 ();
 sg13g2_fill_1 FILLER_48_715 ();
 sg13g2_decap_4 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_816 ();
 sg13g2_decap_8 FILLER_48_823 ();
 sg13g2_decap_8 FILLER_48_830 ();
 sg13g2_decap_8 FILLER_48_837 ();
 sg13g2_decap_8 FILLER_48_844 ();
 sg13g2_decap_8 FILLER_48_851 ();
 sg13g2_decap_8 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_48_865 ();
 sg13g2_decap_8 FILLER_48_872 ();
 sg13g2_decap_8 FILLER_48_879 ();
 sg13g2_decap_8 FILLER_48_886 ();
 sg13g2_decap_8 FILLER_48_893 ();
 sg13g2_decap_8 FILLER_48_900 ();
 sg13g2_decap_8 FILLER_48_907 ();
 sg13g2_decap_8 FILLER_48_914 ();
 sg13g2_decap_8 FILLER_48_921 ();
 sg13g2_decap_8 FILLER_48_928 ();
 sg13g2_decap_8 FILLER_48_935 ();
 sg13g2_decap_8 FILLER_48_942 ();
 sg13g2_decap_8 FILLER_48_949 ();
 sg13g2_decap_8 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_decap_8 FILLER_48_970 ();
 sg13g2_decap_8 FILLER_48_977 ();
 sg13g2_decap_8 FILLER_48_984 ();
 sg13g2_decap_8 FILLER_48_991 ();
 sg13g2_decap_8 FILLER_48_998 ();
 sg13g2_decap_8 FILLER_48_1005 ();
 sg13g2_decap_8 FILLER_48_1012 ();
 sg13g2_decap_8 FILLER_48_1019 ();
 sg13g2_fill_2 FILLER_48_1026 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_decap_8 FILLER_49_114 ();
 sg13g2_decap_8 FILLER_49_121 ();
 sg13g2_decap_8 FILLER_49_128 ();
 sg13g2_decap_8 FILLER_49_143 ();
 sg13g2_decap_8 FILLER_49_150 ();
 sg13g2_decap_8 FILLER_49_157 ();
 sg13g2_decap_8 FILLER_49_164 ();
 sg13g2_decap_8 FILLER_49_171 ();
 sg13g2_decap_8 FILLER_49_178 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_decap_8 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_215 ();
 sg13g2_decap_8 FILLER_49_220 ();
 sg13g2_decap_8 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_234 ();
 sg13g2_decap_8 FILLER_49_241 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_fill_2 FILLER_49_259 ();
 sg13g2_decap_4 FILLER_49_265 ();
 sg13g2_fill_2 FILLER_49_269 ();
 sg13g2_decap_4 FILLER_49_275 ();
 sg13g2_decap_8 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_290 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_decap_8 FILLER_49_302 ();
 sg13g2_decap_8 FILLER_49_309 ();
 sg13g2_decap_4 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_320 ();
 sg13g2_decap_4 FILLER_49_330 ();
 sg13g2_fill_1 FILLER_49_334 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_decap_4 FILLER_49_352 ();
 sg13g2_decap_8 FILLER_49_360 ();
 sg13g2_decap_4 FILLER_49_367 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_8 FILLER_49_404 ();
 sg13g2_decap_8 FILLER_49_411 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_decap_8 FILLER_49_425 ();
 sg13g2_fill_1 FILLER_49_432 ();
 sg13g2_decap_8 FILLER_49_437 ();
 sg13g2_decap_8 FILLER_49_444 ();
 sg13g2_decap_8 FILLER_49_451 ();
 sg13g2_decap_8 FILLER_49_458 ();
 sg13g2_decap_8 FILLER_49_465 ();
 sg13g2_decap_4 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_476 ();
 sg13g2_decap_4 FILLER_49_481 ();
 sg13g2_fill_1 FILLER_49_485 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_4 FILLER_49_497 ();
 sg13g2_fill_1 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_506 ();
 sg13g2_decap_8 FILLER_49_513 ();
 sg13g2_decap_8 FILLER_49_520 ();
 sg13g2_decap_8 FILLER_49_527 ();
 sg13g2_decap_8 FILLER_49_534 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_decap_8 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_decap_8 FILLER_49_569 ();
 sg13g2_decap_8 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_583 ();
 sg13g2_decap_8 FILLER_49_590 ();
 sg13g2_decap_8 FILLER_49_597 ();
 sg13g2_decap_8 FILLER_49_613 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_4 FILLER_49_627 ();
 sg13g2_fill_2 FILLER_49_631 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_fill_2 FILLER_49_649 ();
 sg13g2_fill_2 FILLER_49_674 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_fill_1 FILLER_49_713 ();
 sg13g2_fill_2 FILLER_49_741 ();
 sg13g2_decap_4 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net19;
 assign uio_oe[1] = net20;
 assign uio_oe[2] = net21;
 assign uio_oe[3] = net22;
 assign uio_oe[4] = net23;
 assign uio_oe[5] = net24;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net26;
 assign uio_out[1] = net27;
 assign uio_out[5] = net28;
 assign uio_out[6] = net29;
 assign uio_out[7] = net30;
endmodule
