-- TEROSHDL Documentation:
--! @title Video Timing Generator
--! @author Pascal G. (gfcwfzkm)
--! @version 1.0
--! @date 18.03.2024
--! @brief Generates the video timing signals for a HDMI output.
--!
--! Developed for the BFH oscilloscope project.
--!
--! This module generates the video timing signals for a VGA-timing compatible HDMI output.
--! It is important that the right pixel timing is used in the generic parameters.
--! The module generates the following signals:
--! - disp_active: Active-high signal indicating that the current pixel is within the visible area
--! - disp_x: Current pixel position in the horizontal direction
--! - disp_y: Current pixel position in the vertical direction
--! - frame_end: Strobe signal, active for one cycle when disp_x = H_VISIBLE
--! - line_end: Strobe signal, active for one cycle when disp_x = H_VISIBLE AND disp_y = V_VISIBLE
--! - hdmi_vsync: Active-high signal indicating the vertical sync pulse
--! - hdmi_hsync: Active-high signal indicating the horizontal sync pulse
--! - hdmi_de: Active-high signal indicating the data enable signal
--! 
--! A single, horizontal line is generated by displaying the color data with the hdmi clock, followed
--! by a front porch, sync pulse and back porch, before a new line can be drawn on the screen:
--!
--! ![Single Line Drawing](https://web.mit.edu/6.111/www/s2004/NEWKIT/images/vga_line.png)
--!
--! Many of these lines form the overall image, where the vertical line generation
--! also follows a structure of various lines with the image data, followed by 
--! a front porch, sync pulse and back porch, before a new image can be drawn:
--!
--! ![Vertical Drawing Process](https://web.mit.edu/6.111/www/s2004/NEWKIT/images/vga_frame.png)
--!
--! Ressources:
--! - https://digilent.com/reference/learn/programmable-logic/tutorials/vga-display-congroller/start 
--! - http://martin.hinner.info/vga/vga.html
--! - https://projectf.io/posts/video-timings-vga-720p-1080p/#hd-1280x720-60-hz
--! - https://web.mit.edu/6.111/www/s2004/NEWKIT/vga.shtml

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.log2;
use ieee.math_real.ceil;

entity vtgen is
    generic (
        H_VISIBLE   : positive := 1280; --! Horizontal resolution
        H_FPORCH    : positive := 110;  --! Horizontal Front Porch
        H_SYNC      : positive := 40;   --! Horizontal Sync Pulse
        H_BPORCH    : positive := 220;  --! Horizontal Back Porch

        V_VISIBLE   : positive := 720;  --! Vertical resolution
        V_FPORCH    : positive := 5;    --! Vertical Front Porch
        V_SYNC      : positive := 5;    --! Vertical Sync Pulse
        V_BPORCH    : positive := 20    --! Vertical Back Porch
    );
    port (
        --! Clock speed required to generate the video signal
        clk   : in std_logic;
        --! Ansynchronous, active-high reset
        reset : in std_logic;

        --! Display-Active signal (active-high)
        disp_active : out std_logic;
        --! Currently drawn pixel position. Can be used to control the RGB by an higher architecture
        disp_x      : out unsigned(integer(ceil(log2(real(H_VISIBLE+H_FPORCH+H_SYNC+H_BPORCH))))-1 downto 0);
        --! Currently drawn pixel position. Can be used to control the RGB by an higher architecture
        disp_y      : out unsigned(integer(ceil(log2(real(V_VISIBLE+V_FPORCH+V_SYNC+V_BPORCH))))-1 downto 0);

        --! Frame End signal (active for one cycle)
        frame_end   : out std_logic;
        --! Line End signal (active for one cycle)
        line_end    : out std_logic;

        --! HDMI V-SYNC signal
        hdmi_vsync  : out std_logic;
        --! HDMI H-SYNC signal
        hdmi_hsync  : out std_logic;
        --! HDMI DataEnable Signal
        hdmi_de     : out std_logic
    );
end entity vtgen;

architecture rtl of vtgen is
    -- Constants for the pixel position calculation
    --! Horizontal pixel position drawing end
    constant H_DRAWING_END  : positive := (H_VISIBLE - 1);
    --! Horizontal pixel position sync start
    constant H_SYNC_START   : positive := (H_DRAWING_END + H_FPORCH);
    --! Horizontal pixel position sync end
    constant H_SYNC_END     : positive := (H_SYNC_START + H_SYNC);
    --! Maximum horizontal pixel position
    constant H_MAX : positive := (H_SYNC_END+H_BPORCH);

    --! Vertical pixel position drawing end
    constant V_DRAWING_END  : positive := (V_VISIBLE - 1);
    --! Vertical pixel position sync start
    constant V_SYNC_START   : positive := (V_DRAWING_END + V_FPORCH);
    --! Vertical pixel position sync end
    constant V_SYNC_END     : positive := (V_SYNC_START + V_SYNC);
    --! Maximum vertical pixel position
    constant V_MAX : positive := (V_SYNC_END+V_BPORCH) - 1;

    --! Pixel X position register
    signal disp_x_reg : unsigned(integer(ceil(log2(real(H_MAX))))-1 downto 0);
    --! Pixel Y position register
    signal disp_y_reg : unsigned(integer(ceil(log2(real(V_MAX))))-1 downto 0);
begin
    --! Output of the coordinates
    disp_x <= disp_x_reg;
    disp_y <= disp_y_reg;

    --! Pixel Position Counter
    --! Increments the pixel position registers
    PIXELCNT : process (clk, reset) is begin
        if rising_edge(clk) then
            if reset = '1' then
                disp_x_reg <= (others => '0');
                disp_y_reg <= (others => '0');
            else
                if (disp_x_reg = H_MAX) then
                    disp_x_reg <= (others => '0');
                    if (disp_y_reg = V_MAX) then
                        disp_y_reg <= (others => '0');
                    else
                        disp_y_reg <= disp_y_reg + 1;
                    end if;
                else
                    disp_x_reg <= disp_x_reg + 1;
                end if;
            end if;
        end if;
    end process PIXELCNT;

    --! Sync Signal Generator
    --! Generates the sync signals for the HDMI output
    SYNCGEN : process (disp_x_reg, disp_y_reg) is begin
        hdmi_vsync <= '1';
        hdmi_hsync <= '1';
        hdmi_de <= '0';
        disp_active <= '1';
        line_end <= '0';
        frame_end <= '0';

        if (disp_x_reg >= H_SYNC_START) and (disp_x_reg < H_SYNC_END) then
            hdmi_hsync <= '0';
        end if;

        if (disp_y_reg >= V_SYNC_START) and (disp_y_reg < V_SYNC_END) then
            hdmi_vsync <= '0';
        end if;

        if (disp_x_reg <= H_DRAWING_END) and (disp_y_reg <= V_DRAWING_END) then
            hdmi_de <= '1';
        end if;

        if (disp_x_reg > H_DRAWING_END) or (disp_y_reg > V_DRAWING_END) then
            disp_active <= '0';
        end if;

        if disp_x_reg = H_VISIBLE then
            if disp_y_reg = V_VISIBLE then
                frame_end <= '1';
            else
                line_end <= '1';
            end if;
        end if;

    end process SYNCGEN;

end architecture;